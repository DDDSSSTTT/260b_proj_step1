##
## LEF for PtnCells ;
## created by Innovus v19.17-s077_1 on Tue Mar 14 18:57:57 2023
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fullchip
  CLASS BLOCK ;
  SIZE 470.000000 BY 466.400000 ;
  FOREIGN fullchip 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 24.950000 0.520000 25.050000 ;
    END
  END clk
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 429.950000 0.520000 430.050000 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 424.950000 0.520000 425.050000 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 419.950000 0.520000 420.050000 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 414.950000 0.520000 415.050000 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 409.950000 0.520000 410.050000 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 404.950000 0.520000 405.050000 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 399.950000 0.520000 400.050000 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 394.950000 0.520000 395.050000 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 389.950000 0.520000 390.050000 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 384.950000 0.520000 385.050000 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 379.950000 0.520000 380.050000 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 374.950000 0.520000 375.050000 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 369.950000 0.520000 370.050000 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 364.950000 0.520000 365.050000 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 359.950000 0.520000 360.050000 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 354.950000 0.520000 355.050000 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 349.950000 0.520000 350.050000 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 344.950000 0.520000 345.050000 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 339.950000 0.520000 340.050000 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 334.950000 0.520000 335.050000 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 329.950000 0.520000 330.050000 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 324.950000 0.520000 325.050000 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 319.950000 0.520000 320.050000 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 314.950000 0.520000 315.050000 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 309.950000 0.520000 310.050000 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 304.950000 0.520000 305.050000 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 299.950000 0.520000 300.050000 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 294.950000 0.520000 295.050000 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 289.950000 0.520000 290.050000 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 284.950000 0.520000 285.050000 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 279.950000 0.520000 280.050000 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 274.950000 0.520000 275.050000 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 269.950000 0.520000 270.050000 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 264.950000 0.520000 265.050000 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 259.950000 0.520000 260.050000 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 254.950000 0.520000 255.050000 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 249.950000 0.520000 250.050000 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 244.950000 0.520000 245.050000 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 239.950000 0.520000 240.050000 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 234.950000 0.520000 235.050000 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 229.950000 0.520000 230.050000 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 224.950000 0.520000 225.050000 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 219.950000 0.520000 220.050000 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 214.950000 0.520000 215.050000 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 209.950000 0.520000 210.050000 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 204.950000 0.520000 205.050000 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 199.950000 0.520000 200.050000 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 194.950000 0.520000 195.050000 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 189.950000 0.520000 190.050000 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 184.950000 0.520000 185.050000 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 179.950000 0.520000 180.050000 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 174.950000 0.520000 175.050000 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 169.950000 0.520000 170.050000 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 164.950000 0.520000 165.050000 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 159.950000 0.520000 160.050000 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 154.950000 0.520000 155.050000 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 149.950000 0.520000 150.050000 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 144.950000 0.520000 145.050000 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 139.950000 0.520000 140.050000 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 134.950000 0.520000 135.050000 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 129.950000 0.520000 130.050000 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 124.950000 0.520000 125.050000 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 119.950000 0.520000 120.050000 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 114.950000 0.520000 115.050000 ;
    END
  END mem_in[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 109.950000 0.520000 110.050000 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 104.950000 0.520000 105.050000 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 99.950000 0.520000 100.050000 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 94.950000 0.520000 95.050000 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 89.950000 0.520000 90.050000 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 84.950000 0.520000 85.050000 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 79.950000 0.520000 80.050000 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 74.950000 0.520000 75.050000 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 69.950000 0.520000 70.050000 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 64.950000 0.520000 65.050000 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 59.950000 0.520000 60.050000 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 54.950000 0.520000 55.050000 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 49.950000 0.520000 50.050000 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 44.950000 0.520000 45.050000 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 39.950000 0.520000 40.050000 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 34.950000 0.520000 35.050000 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 29.950000 0.520000 30.050000 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 434.950000 0.520000 435.050000 ;
    END
  END reset
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.850000 0.000000 159.950000 0.520000 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.850000 0.000000 162.950000 0.520000 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.850000 0.000000 165.950000 0.520000 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.850000 0.000000 168.950000 0.520000 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.850000 0.000000 171.950000 0.520000 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 174.850000 0.000000 174.950000 0.520000 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.850000 0.000000 177.950000 0.520000 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 180.850000 0.000000 180.950000 0.520000 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.850000 0.000000 183.950000 0.520000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.850000 0.000000 186.950000 0.520000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 189.850000 0.000000 189.950000 0.520000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 192.850000 0.000000 192.950000 0.520000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 195.850000 0.000000 195.950000 0.520000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 198.850000 0.000000 198.950000 0.520000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 201.850000 0.000000 201.950000 0.520000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.850000 0.000000 204.950000 0.520000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.850000 0.000000 207.950000 0.520000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 210.850000 0.000000 210.950000 0.520000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 213.850000 0.000000 213.950000 0.520000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.850000 0.000000 216.950000 0.520000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.850000 0.000000 219.950000 0.520000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 222.850000 0.000000 222.950000 0.520000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 225.850000 0.000000 225.950000 0.520000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 228.850000 0.000000 228.950000 0.520000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 231.850000 0.000000 231.950000 0.520000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 234.850000 0.000000 234.950000 0.520000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 237.850000 0.000000 237.950000 0.520000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 240.850000 0.000000 240.950000 0.520000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 243.850000 0.000000 243.950000 0.520000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 246.850000 0.000000 246.950000 0.520000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 249.850000 0.000000 249.950000 0.520000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 252.850000 0.000000 252.950000 0.520000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 255.850000 0.000000 255.950000 0.520000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 258.850000 0.000000 258.950000 0.520000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 261.850000 0.000000 261.950000 0.520000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 264.850000 0.000000 264.950000 0.520000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 267.850000 0.000000 267.950000 0.520000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 270.850000 0.000000 270.950000 0.520000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 273.850000 0.000000 273.950000 0.520000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 276.850000 0.000000 276.950000 0.520000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 279.850000 0.000000 279.950000 0.520000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 282.850000 0.000000 282.950000 0.520000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 285.850000 0.000000 285.950000 0.520000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 288.850000 0.000000 288.950000 0.520000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 291.850000 0.000000 291.950000 0.520000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 294.850000 0.000000 294.950000 0.520000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 297.850000 0.000000 297.950000 0.520000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 300.850000 0.000000 300.950000 0.520000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 303.850000 0.000000 303.950000 0.520000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 306.850000 0.000000 306.950000 0.520000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 309.850000 0.000000 309.950000 0.520000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 312.850000 0.000000 312.950000 0.520000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 315.850000 0.000000 315.950000 0.520000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 318.850000 0.000000 318.950000 0.520000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 321.850000 0.000000 321.950000 0.520000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 324.850000 0.000000 324.950000 0.520000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 327.850000 0.000000 327.950000 0.520000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 330.850000 0.000000 330.950000 0.520000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 333.850000 0.000000 333.950000 0.520000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 336.850000 0.000000 336.950000 0.520000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.850000 0.000000 339.950000 0.520000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 342.850000 0.000000 342.950000 0.520000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 345.850000 0.000000 345.950000 0.520000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 348.850000 0.000000 348.950000 0.520000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 351.850000 0.000000 351.950000 0.520000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 354.850000 0.000000 354.950000 0.520000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 357.850000 0.000000 357.950000 0.520000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 360.850000 0.000000 360.950000 0.520000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 363.850000 0.000000 363.950000 0.520000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 366.850000 0.000000 366.950000 0.520000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 369.850000 0.000000 369.950000 0.520000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 372.850000 0.000000 372.950000 0.520000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 375.850000 0.000000 375.950000 0.520000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 378.850000 0.000000 378.950000 0.520000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 381.850000 0.000000 381.950000 0.520000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 384.850000 0.000000 384.950000 0.520000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 387.850000 0.000000 387.950000 0.520000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 390.850000 0.000000 390.950000 0.520000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 393.850000 0.000000 393.950000 0.520000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 396.850000 0.000000 396.950000 0.520000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 399.850000 0.000000 399.950000 0.520000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 402.850000 0.000000 402.950000 0.520000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 405.850000 0.000000 405.950000 0.520000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 408.850000 0.000000 408.950000 0.520000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 411.850000 0.000000 411.950000 0.520000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 414.850000 0.000000 414.950000 0.520000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 417.850000 0.000000 417.950000 0.520000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 420.850000 0.000000 420.950000 0.520000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 423.850000 0.000000 423.950000 0.520000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 426.850000 0.000000 426.950000 0.520000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 429.850000 0.000000 429.950000 0.520000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 432.850000 0.000000 432.950000 0.520000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 435.850000 0.000000 435.950000 0.520000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 438.850000 0.000000 438.950000 0.520000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 441.850000 0.000000 441.950000 0.520000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 444.850000 0.000000 444.950000 0.520000 ;
    END
  END out[0]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.850000 0.000000 111.950000 0.520000 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.850000 0.000000 114.950000 0.520000 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.850000 0.000000 117.950000 0.520000 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.850000 0.000000 120.950000 0.520000 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.850000 0.000000 123.950000 0.520000 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.850000 0.000000 126.950000 0.520000 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.850000 0.000000 129.950000 0.520000 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.850000 0.000000 132.950000 0.520000 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.850000 0.000000 135.950000 0.520000 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.850000 0.000000 138.950000 0.520000 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.850000 0.000000 141.950000 0.520000 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.850000 0.000000 144.950000 0.520000 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.850000 0.000000 147.950000 0.520000 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.850000 0.000000 150.950000 0.520000 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.850000 0.000000 153.950000 0.520000 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.850000 0.000000 156.950000 0.520000 ;
    END
  END sum_out[0]
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 470.000000 466.400000 ;
    LAYER M2 ;
      RECT 0.000000 0.640000 470.000000 466.400000 ;
      RECT 445.050000 0.000000 470.000000 0.640000 ;
      RECT 442.050000 0.000000 444.750000 0.640000 ;
      RECT 439.050000 0.000000 441.750000 0.640000 ;
      RECT 436.050000 0.000000 438.750000 0.640000 ;
      RECT 433.050000 0.000000 435.750000 0.640000 ;
      RECT 430.050000 0.000000 432.750000 0.640000 ;
      RECT 427.050000 0.000000 429.750000 0.640000 ;
      RECT 424.050000 0.000000 426.750000 0.640000 ;
      RECT 421.050000 0.000000 423.750000 0.640000 ;
      RECT 418.050000 0.000000 420.750000 0.640000 ;
      RECT 415.050000 0.000000 417.750000 0.640000 ;
      RECT 412.050000 0.000000 414.750000 0.640000 ;
      RECT 409.050000 0.000000 411.750000 0.640000 ;
      RECT 406.050000 0.000000 408.750000 0.640000 ;
      RECT 403.050000 0.000000 405.750000 0.640000 ;
      RECT 400.050000 0.000000 402.750000 0.640000 ;
      RECT 397.050000 0.000000 399.750000 0.640000 ;
      RECT 394.050000 0.000000 396.750000 0.640000 ;
      RECT 391.050000 0.000000 393.750000 0.640000 ;
      RECT 388.050000 0.000000 390.750000 0.640000 ;
      RECT 385.050000 0.000000 387.750000 0.640000 ;
      RECT 382.050000 0.000000 384.750000 0.640000 ;
      RECT 379.050000 0.000000 381.750000 0.640000 ;
      RECT 376.050000 0.000000 378.750000 0.640000 ;
      RECT 373.050000 0.000000 375.750000 0.640000 ;
      RECT 370.050000 0.000000 372.750000 0.640000 ;
      RECT 367.050000 0.000000 369.750000 0.640000 ;
      RECT 364.050000 0.000000 366.750000 0.640000 ;
      RECT 361.050000 0.000000 363.750000 0.640000 ;
      RECT 358.050000 0.000000 360.750000 0.640000 ;
      RECT 355.050000 0.000000 357.750000 0.640000 ;
      RECT 352.050000 0.000000 354.750000 0.640000 ;
      RECT 349.050000 0.000000 351.750000 0.640000 ;
      RECT 346.050000 0.000000 348.750000 0.640000 ;
      RECT 343.050000 0.000000 345.750000 0.640000 ;
      RECT 340.050000 0.000000 342.750000 0.640000 ;
      RECT 337.050000 0.000000 339.750000 0.640000 ;
      RECT 334.050000 0.000000 336.750000 0.640000 ;
      RECT 331.050000 0.000000 333.750000 0.640000 ;
      RECT 328.050000 0.000000 330.750000 0.640000 ;
      RECT 325.050000 0.000000 327.750000 0.640000 ;
      RECT 322.050000 0.000000 324.750000 0.640000 ;
      RECT 319.050000 0.000000 321.750000 0.640000 ;
      RECT 316.050000 0.000000 318.750000 0.640000 ;
      RECT 313.050000 0.000000 315.750000 0.640000 ;
      RECT 310.050000 0.000000 312.750000 0.640000 ;
      RECT 307.050000 0.000000 309.750000 0.640000 ;
      RECT 304.050000 0.000000 306.750000 0.640000 ;
      RECT 301.050000 0.000000 303.750000 0.640000 ;
      RECT 298.050000 0.000000 300.750000 0.640000 ;
      RECT 295.050000 0.000000 297.750000 0.640000 ;
      RECT 292.050000 0.000000 294.750000 0.640000 ;
      RECT 289.050000 0.000000 291.750000 0.640000 ;
      RECT 286.050000 0.000000 288.750000 0.640000 ;
      RECT 283.050000 0.000000 285.750000 0.640000 ;
      RECT 280.050000 0.000000 282.750000 0.640000 ;
      RECT 277.050000 0.000000 279.750000 0.640000 ;
      RECT 274.050000 0.000000 276.750000 0.640000 ;
      RECT 271.050000 0.000000 273.750000 0.640000 ;
      RECT 268.050000 0.000000 270.750000 0.640000 ;
      RECT 265.050000 0.000000 267.750000 0.640000 ;
      RECT 262.050000 0.000000 264.750000 0.640000 ;
      RECT 259.050000 0.000000 261.750000 0.640000 ;
      RECT 256.050000 0.000000 258.750000 0.640000 ;
      RECT 253.050000 0.000000 255.750000 0.640000 ;
      RECT 250.050000 0.000000 252.750000 0.640000 ;
      RECT 247.050000 0.000000 249.750000 0.640000 ;
      RECT 244.050000 0.000000 246.750000 0.640000 ;
      RECT 241.050000 0.000000 243.750000 0.640000 ;
      RECT 238.050000 0.000000 240.750000 0.640000 ;
      RECT 235.050000 0.000000 237.750000 0.640000 ;
      RECT 232.050000 0.000000 234.750000 0.640000 ;
      RECT 229.050000 0.000000 231.750000 0.640000 ;
      RECT 226.050000 0.000000 228.750000 0.640000 ;
      RECT 223.050000 0.000000 225.750000 0.640000 ;
      RECT 220.050000 0.000000 222.750000 0.640000 ;
      RECT 217.050000 0.000000 219.750000 0.640000 ;
      RECT 214.050000 0.000000 216.750000 0.640000 ;
      RECT 211.050000 0.000000 213.750000 0.640000 ;
      RECT 208.050000 0.000000 210.750000 0.640000 ;
      RECT 205.050000 0.000000 207.750000 0.640000 ;
      RECT 202.050000 0.000000 204.750000 0.640000 ;
      RECT 199.050000 0.000000 201.750000 0.640000 ;
      RECT 196.050000 0.000000 198.750000 0.640000 ;
      RECT 193.050000 0.000000 195.750000 0.640000 ;
      RECT 190.050000 0.000000 192.750000 0.640000 ;
      RECT 187.050000 0.000000 189.750000 0.640000 ;
      RECT 184.050000 0.000000 186.750000 0.640000 ;
      RECT 181.050000 0.000000 183.750000 0.640000 ;
      RECT 178.050000 0.000000 180.750000 0.640000 ;
      RECT 175.050000 0.000000 177.750000 0.640000 ;
      RECT 172.050000 0.000000 174.750000 0.640000 ;
      RECT 169.050000 0.000000 171.750000 0.640000 ;
      RECT 166.050000 0.000000 168.750000 0.640000 ;
      RECT 163.050000 0.000000 165.750000 0.640000 ;
      RECT 160.050000 0.000000 162.750000 0.640000 ;
      RECT 157.050000 0.000000 159.750000 0.640000 ;
      RECT 154.050000 0.000000 156.750000 0.640000 ;
      RECT 151.050000 0.000000 153.750000 0.640000 ;
      RECT 148.050000 0.000000 150.750000 0.640000 ;
      RECT 145.050000 0.000000 147.750000 0.640000 ;
      RECT 142.050000 0.000000 144.750000 0.640000 ;
      RECT 139.050000 0.000000 141.750000 0.640000 ;
      RECT 136.050000 0.000000 138.750000 0.640000 ;
      RECT 133.050000 0.000000 135.750000 0.640000 ;
      RECT 130.050000 0.000000 132.750000 0.640000 ;
      RECT 127.050000 0.000000 129.750000 0.640000 ;
      RECT 124.050000 0.000000 126.750000 0.640000 ;
      RECT 121.050000 0.000000 123.750000 0.640000 ;
      RECT 118.050000 0.000000 120.750000 0.640000 ;
      RECT 115.050000 0.000000 117.750000 0.640000 ;
      RECT 112.050000 0.000000 114.750000 0.640000 ;
      RECT 0.000000 0.000000 111.750000 0.640000 ;
    LAYER M3 ;
      RECT 0.000000 435.150000 470.000000 466.400000 ;
      RECT 0.640000 434.850000 470.000000 435.150000 ;
      RECT 0.000000 430.150000 470.000000 434.850000 ;
      RECT 0.640000 429.850000 470.000000 430.150000 ;
      RECT 0.000000 425.150000 470.000000 429.850000 ;
      RECT 0.640000 424.850000 470.000000 425.150000 ;
      RECT 0.000000 420.150000 470.000000 424.850000 ;
      RECT 0.640000 419.850000 470.000000 420.150000 ;
      RECT 0.000000 415.150000 470.000000 419.850000 ;
      RECT 0.640000 414.850000 470.000000 415.150000 ;
      RECT 0.000000 410.150000 470.000000 414.850000 ;
      RECT 0.640000 409.850000 470.000000 410.150000 ;
      RECT 0.000000 405.150000 470.000000 409.850000 ;
      RECT 0.640000 404.850000 470.000000 405.150000 ;
      RECT 0.000000 400.150000 470.000000 404.850000 ;
      RECT 0.640000 399.850000 470.000000 400.150000 ;
      RECT 0.000000 395.150000 470.000000 399.850000 ;
      RECT 0.640000 394.850000 470.000000 395.150000 ;
      RECT 0.000000 390.150000 470.000000 394.850000 ;
      RECT 0.640000 389.850000 470.000000 390.150000 ;
      RECT 0.000000 385.150000 470.000000 389.850000 ;
      RECT 0.640000 384.850000 470.000000 385.150000 ;
      RECT 0.000000 380.150000 470.000000 384.850000 ;
      RECT 0.640000 379.850000 470.000000 380.150000 ;
      RECT 0.000000 375.150000 470.000000 379.850000 ;
      RECT 0.640000 374.850000 470.000000 375.150000 ;
      RECT 0.000000 370.150000 470.000000 374.850000 ;
      RECT 0.640000 369.850000 470.000000 370.150000 ;
      RECT 0.000000 365.150000 470.000000 369.850000 ;
      RECT 0.640000 364.850000 470.000000 365.150000 ;
      RECT 0.000000 360.150000 470.000000 364.850000 ;
      RECT 0.640000 359.850000 470.000000 360.150000 ;
      RECT 0.000000 355.150000 470.000000 359.850000 ;
      RECT 0.640000 354.850000 470.000000 355.150000 ;
      RECT 0.000000 350.150000 470.000000 354.850000 ;
      RECT 0.640000 349.850000 470.000000 350.150000 ;
      RECT 0.000000 345.150000 470.000000 349.850000 ;
      RECT 0.640000 344.850000 470.000000 345.150000 ;
      RECT 0.000000 340.150000 470.000000 344.850000 ;
      RECT 0.640000 339.850000 470.000000 340.150000 ;
      RECT 0.000000 335.150000 470.000000 339.850000 ;
      RECT 0.640000 334.850000 470.000000 335.150000 ;
      RECT 0.000000 330.150000 470.000000 334.850000 ;
      RECT 0.640000 329.850000 470.000000 330.150000 ;
      RECT 0.000000 325.150000 470.000000 329.850000 ;
      RECT 0.640000 324.850000 470.000000 325.150000 ;
      RECT 0.000000 320.150000 470.000000 324.850000 ;
      RECT 0.640000 319.850000 470.000000 320.150000 ;
      RECT 0.000000 315.150000 470.000000 319.850000 ;
      RECT 0.640000 314.850000 470.000000 315.150000 ;
      RECT 0.000000 310.150000 470.000000 314.850000 ;
      RECT 0.640000 309.850000 470.000000 310.150000 ;
      RECT 0.000000 305.150000 470.000000 309.850000 ;
      RECT 0.640000 304.850000 470.000000 305.150000 ;
      RECT 0.000000 300.150000 470.000000 304.850000 ;
      RECT 0.640000 299.850000 470.000000 300.150000 ;
      RECT 0.000000 295.150000 470.000000 299.850000 ;
      RECT 0.640000 294.850000 470.000000 295.150000 ;
      RECT 0.000000 290.150000 470.000000 294.850000 ;
      RECT 0.640000 289.850000 470.000000 290.150000 ;
      RECT 0.000000 285.150000 470.000000 289.850000 ;
      RECT 0.640000 284.850000 470.000000 285.150000 ;
      RECT 0.000000 280.150000 470.000000 284.850000 ;
      RECT 0.640000 279.850000 470.000000 280.150000 ;
      RECT 0.000000 275.150000 470.000000 279.850000 ;
      RECT 0.640000 274.850000 470.000000 275.150000 ;
      RECT 0.000000 270.150000 470.000000 274.850000 ;
      RECT 0.640000 269.850000 470.000000 270.150000 ;
      RECT 0.000000 265.150000 470.000000 269.850000 ;
      RECT 0.640000 264.850000 470.000000 265.150000 ;
      RECT 0.000000 260.150000 470.000000 264.850000 ;
      RECT 0.640000 259.850000 470.000000 260.150000 ;
      RECT 0.000000 255.150000 470.000000 259.850000 ;
      RECT 0.640000 254.850000 470.000000 255.150000 ;
      RECT 0.000000 250.150000 470.000000 254.850000 ;
      RECT 0.640000 249.850000 470.000000 250.150000 ;
      RECT 0.000000 245.150000 470.000000 249.850000 ;
      RECT 0.640000 244.850000 470.000000 245.150000 ;
      RECT 0.000000 240.150000 470.000000 244.850000 ;
      RECT 0.640000 239.850000 470.000000 240.150000 ;
      RECT 0.000000 235.150000 470.000000 239.850000 ;
      RECT 0.640000 234.850000 470.000000 235.150000 ;
      RECT 0.000000 230.150000 470.000000 234.850000 ;
      RECT 0.640000 229.850000 470.000000 230.150000 ;
      RECT 0.000000 225.150000 470.000000 229.850000 ;
      RECT 0.640000 224.850000 470.000000 225.150000 ;
      RECT 0.000000 220.150000 470.000000 224.850000 ;
      RECT 0.640000 219.850000 470.000000 220.150000 ;
      RECT 0.000000 215.150000 470.000000 219.850000 ;
      RECT 0.640000 214.850000 470.000000 215.150000 ;
      RECT 0.000000 210.150000 470.000000 214.850000 ;
      RECT 0.640000 209.850000 470.000000 210.150000 ;
      RECT 0.000000 205.150000 470.000000 209.850000 ;
      RECT 0.640000 204.850000 470.000000 205.150000 ;
      RECT 0.000000 200.150000 470.000000 204.850000 ;
      RECT 0.640000 199.850000 470.000000 200.150000 ;
      RECT 0.000000 195.150000 470.000000 199.850000 ;
      RECT 0.640000 194.850000 470.000000 195.150000 ;
      RECT 0.000000 190.150000 470.000000 194.850000 ;
      RECT 0.640000 189.850000 470.000000 190.150000 ;
      RECT 0.000000 185.150000 470.000000 189.850000 ;
      RECT 0.640000 184.850000 470.000000 185.150000 ;
      RECT 0.000000 180.150000 470.000000 184.850000 ;
      RECT 0.640000 179.850000 470.000000 180.150000 ;
      RECT 0.000000 175.150000 470.000000 179.850000 ;
      RECT 0.640000 174.850000 470.000000 175.150000 ;
      RECT 0.000000 170.150000 470.000000 174.850000 ;
      RECT 0.640000 169.850000 470.000000 170.150000 ;
      RECT 0.000000 165.150000 470.000000 169.850000 ;
      RECT 0.640000 164.850000 470.000000 165.150000 ;
      RECT 0.000000 160.150000 470.000000 164.850000 ;
      RECT 0.640000 159.850000 470.000000 160.150000 ;
      RECT 0.000000 155.150000 470.000000 159.850000 ;
      RECT 0.640000 154.850000 470.000000 155.150000 ;
      RECT 0.000000 150.150000 470.000000 154.850000 ;
      RECT 0.640000 149.850000 470.000000 150.150000 ;
      RECT 0.000000 145.150000 470.000000 149.850000 ;
      RECT 0.640000 144.850000 470.000000 145.150000 ;
      RECT 0.000000 140.150000 470.000000 144.850000 ;
      RECT 0.640000 139.850000 470.000000 140.150000 ;
      RECT 0.000000 135.150000 470.000000 139.850000 ;
      RECT 0.640000 134.850000 470.000000 135.150000 ;
      RECT 0.000000 130.150000 470.000000 134.850000 ;
      RECT 0.640000 129.850000 470.000000 130.150000 ;
      RECT 0.000000 125.150000 470.000000 129.850000 ;
      RECT 0.640000 124.850000 470.000000 125.150000 ;
      RECT 0.000000 120.150000 470.000000 124.850000 ;
      RECT 0.640000 119.850000 470.000000 120.150000 ;
      RECT 0.000000 115.150000 470.000000 119.850000 ;
      RECT 0.640000 114.850000 470.000000 115.150000 ;
      RECT 0.000000 110.150000 470.000000 114.850000 ;
      RECT 0.640000 109.850000 470.000000 110.150000 ;
      RECT 0.000000 105.150000 470.000000 109.850000 ;
      RECT 0.640000 104.850000 470.000000 105.150000 ;
      RECT 0.000000 100.150000 470.000000 104.850000 ;
      RECT 0.640000 99.850000 470.000000 100.150000 ;
      RECT 0.000000 95.150000 470.000000 99.850000 ;
      RECT 0.640000 94.850000 470.000000 95.150000 ;
      RECT 0.000000 90.150000 470.000000 94.850000 ;
      RECT 0.640000 89.850000 470.000000 90.150000 ;
      RECT 0.000000 85.150000 470.000000 89.850000 ;
      RECT 0.640000 84.850000 470.000000 85.150000 ;
      RECT 0.000000 80.150000 470.000000 84.850000 ;
      RECT 0.640000 79.850000 470.000000 80.150000 ;
      RECT 0.000000 75.150000 470.000000 79.850000 ;
      RECT 0.640000 74.850000 470.000000 75.150000 ;
      RECT 0.000000 70.150000 470.000000 74.850000 ;
      RECT 0.640000 69.850000 470.000000 70.150000 ;
      RECT 0.000000 65.150000 470.000000 69.850000 ;
      RECT 0.640000 64.850000 470.000000 65.150000 ;
      RECT 0.000000 60.150000 470.000000 64.850000 ;
      RECT 0.640000 59.850000 470.000000 60.150000 ;
      RECT 0.000000 55.150000 470.000000 59.850000 ;
      RECT 0.640000 54.850000 470.000000 55.150000 ;
      RECT 0.000000 50.150000 470.000000 54.850000 ;
      RECT 0.640000 49.850000 470.000000 50.150000 ;
      RECT 0.000000 45.150000 470.000000 49.850000 ;
      RECT 0.640000 44.850000 470.000000 45.150000 ;
      RECT 0.000000 40.150000 470.000000 44.850000 ;
      RECT 0.640000 39.850000 470.000000 40.150000 ;
      RECT 0.000000 35.150000 470.000000 39.850000 ;
      RECT 0.640000 34.850000 470.000000 35.150000 ;
      RECT 0.000000 30.150000 470.000000 34.850000 ;
      RECT 0.640000 29.850000 470.000000 30.150000 ;
      RECT 0.000000 25.150000 470.000000 29.850000 ;
      RECT 0.640000 24.850000 470.000000 25.150000 ;
      RECT 0.000000 0.000000 470.000000 24.850000 ;
    LAYER M4 ;
      RECT 0.000000 0.000000 470.000000 466.400000 ;
    LAYER M5 ;
      RECT 0.000000 0.000000 470.000000 466.400000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 470.000000 466.400000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 470.000000 466.400000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 470.000000 466.400000 ;
  END
END fullchip

END LIBRARY
