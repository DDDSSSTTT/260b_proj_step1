##
## LEF for PtnCells ;
## created by Innovus v19.17-s077_1 on Mon Feb 20 13:59:36 2023
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO add
  CLASS BLOCK ;
  SIZE 40.800000 BY 38.000000 ;
  FOREIGN add 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.000000 9.155000 0.470000 9.245000 ;
    END
  END clk
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 40.330000 15.155000 40.800000 15.245000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 40.330000 16.755000 40.800000 16.845000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 40.330000 18.355000 40.800000 18.445000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 40.330000 19.955000 40.800000 20.045000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 40.330000 21.555000 40.800000 21.645000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 40.330000 23.155000 40.800000 23.245000 ;
    END
  END out[0]
  PIN x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.000000 15.555000 0.470000 15.645000 ;
    END
  END x[3]
  PIN x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.000000 13.955000 0.470000 14.045000 ;
    END
  END x[2]
  PIN x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.000000 12.355000 0.470000 12.445000 ;
    END
  END x[1]
  PIN x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.000000 10.755000 0.470000 10.845000 ;
    END
  END x[0]
  PIN y[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.000000 21.955000 0.470000 22.045000 ;
    END
  END y[3]
  PIN y[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.000000 20.355000 0.470000 20.445000 ;
    END
  END y[2]
  PIN y[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.000000 18.755000 0.470000 18.845000 ;
    END
  END y[1]
  PIN y[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.000000 17.155000 0.470000 17.245000 ;
    END
  END y[0]
  PIN z[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.000000 28.355000 0.470000 28.445000 ;
    END
  END z[3]
  PIN z[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.000000 26.755000 0.470000 26.845000 ;
    END
  END z[2]
  PIN z[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.000000 25.155000 0.470000 25.245000 ;
    END
  END z[1]
  PIN z[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.000000 23.555000 0.470000 23.645000 ;
    END
  END z[0]
  OBS
    LAYER M1 ;
      RECT 0.000000 28.535000 40.800000 38.000000 ;
      RECT 0.580000 28.265000 40.800000 28.535000 ;
      RECT 0.000000 26.935000 40.800000 28.265000 ;
      RECT 0.580000 26.665000 40.800000 26.935000 ;
      RECT 0.000000 25.335000 40.800000 26.665000 ;
      RECT 0.580000 25.065000 40.800000 25.335000 ;
      RECT 0.000000 23.735000 40.800000 25.065000 ;
      RECT 0.580000 23.465000 40.800000 23.735000 ;
      RECT 0.000000 23.335000 40.800000 23.465000 ;
      RECT 0.000000 23.065000 40.220000 23.335000 ;
      RECT 0.000000 22.135000 40.800000 23.065000 ;
      RECT 0.580000 21.865000 40.800000 22.135000 ;
      RECT 0.000000 21.735000 40.800000 21.865000 ;
      RECT 0.000000 21.465000 40.220000 21.735000 ;
      RECT 0.000000 20.535000 40.800000 21.465000 ;
      RECT 0.580000 20.265000 40.800000 20.535000 ;
      RECT 0.000000 20.135000 40.800000 20.265000 ;
      RECT 0.000000 19.865000 40.220000 20.135000 ;
      RECT 0.000000 18.935000 40.800000 19.865000 ;
      RECT 0.580000 18.665000 40.800000 18.935000 ;
      RECT 0.000000 18.535000 40.800000 18.665000 ;
      RECT 0.000000 18.265000 40.220000 18.535000 ;
      RECT 0.000000 17.335000 40.800000 18.265000 ;
      RECT 0.580000 17.065000 40.800000 17.335000 ;
      RECT 0.000000 16.935000 40.800000 17.065000 ;
      RECT 0.000000 16.665000 40.220000 16.935000 ;
      RECT 0.000000 15.735000 40.800000 16.665000 ;
      RECT 0.580000 15.465000 40.800000 15.735000 ;
      RECT 0.000000 15.335000 40.800000 15.465000 ;
      RECT 0.000000 15.065000 40.220000 15.335000 ;
      RECT 0.000000 14.135000 40.800000 15.065000 ;
      RECT 0.580000 13.865000 40.800000 14.135000 ;
      RECT 0.000000 12.535000 40.800000 13.865000 ;
      RECT 0.580000 12.265000 40.800000 12.535000 ;
      RECT 0.000000 10.935000 40.800000 12.265000 ;
      RECT 0.580000 10.665000 40.800000 10.935000 ;
      RECT 0.000000 9.335000 40.800000 10.665000 ;
      RECT 0.580000 9.065000 40.800000 9.335000 ;
      RECT 0.000000 0.000000 40.800000 9.065000 ;
    LAYER M2 ;
      RECT 0.000000 0.000000 40.800000 38.000000 ;
    LAYER M3 ;
      RECT 0.000000 0.000000 40.800000 38.000000 ;
    LAYER M4 ;
      RECT 0.000000 0.000000 40.800000 38.000000 ;
    LAYER M5 ;
      RECT 0.000000 0.000000 40.800000 38.000000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 40.800000 38.000000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 40.800000 38.000000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 40.800000 38.000000 ;
  END
END add

END LIBRARY
