##
## LEF for PtnCells ;
## created by Innovus v19.17-s077_1 on Mon Mar 13 00:14:43 2023
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fullchip
  CLASS BLOCK ;
  SIZE 693.200000 BY 689.600000 ;
  FOREIGN fullchip 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 24.950000 0.520000 25.050000 ;
    END
  END clk
  PIN mem_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 314.950000 0.520000 315.050000 ;
    END
  END mem_in[127]
  PIN mem_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 312.950000 0.520000 313.050000 ;
    END
  END mem_in[126]
  PIN mem_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 310.950000 0.520000 311.050000 ;
    END
  END mem_in[125]
  PIN mem_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 308.950000 0.520000 309.050000 ;
    END
  END mem_in[124]
  PIN mem_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 306.950000 0.520000 307.050000 ;
    END
  END mem_in[123]
  PIN mem_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 304.950000 0.520000 305.050000 ;
    END
  END mem_in[122]
  PIN mem_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 302.950000 0.520000 303.050000 ;
    END
  END mem_in[121]
  PIN mem_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 300.950000 0.520000 301.050000 ;
    END
  END mem_in[120]
  PIN mem_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 298.950000 0.520000 299.050000 ;
    END
  END mem_in[119]
  PIN mem_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 296.950000 0.520000 297.050000 ;
    END
  END mem_in[118]
  PIN mem_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 294.950000 0.520000 295.050000 ;
    END
  END mem_in[117]
  PIN mem_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 292.950000 0.520000 293.050000 ;
    END
  END mem_in[116]
  PIN mem_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 290.950000 0.520000 291.050000 ;
    END
  END mem_in[115]
  PIN mem_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 288.950000 0.520000 289.050000 ;
    END
  END mem_in[114]
  PIN mem_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 286.950000 0.520000 287.050000 ;
    END
  END mem_in[113]
  PIN mem_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 284.950000 0.520000 285.050000 ;
    END
  END mem_in[112]
  PIN mem_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 282.950000 0.520000 283.050000 ;
    END
  END mem_in[111]
  PIN mem_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 280.950000 0.520000 281.050000 ;
    END
  END mem_in[110]
  PIN mem_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 278.950000 0.520000 279.050000 ;
    END
  END mem_in[109]
  PIN mem_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 276.950000 0.520000 277.050000 ;
    END
  END mem_in[108]
  PIN mem_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 274.950000 0.520000 275.050000 ;
    END
  END mem_in[107]
  PIN mem_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 272.950000 0.520000 273.050000 ;
    END
  END mem_in[106]
  PIN mem_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 270.950000 0.520000 271.050000 ;
    END
  END mem_in[105]
  PIN mem_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 268.950000 0.520000 269.050000 ;
    END
  END mem_in[104]
  PIN mem_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 266.950000 0.520000 267.050000 ;
    END
  END mem_in[103]
  PIN mem_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 264.950000 0.520000 265.050000 ;
    END
  END mem_in[102]
  PIN mem_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 262.950000 0.520000 263.050000 ;
    END
  END mem_in[101]
  PIN mem_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 260.950000 0.520000 261.050000 ;
    END
  END mem_in[100]
  PIN mem_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 258.950000 0.520000 259.050000 ;
    END
  END mem_in[99]
  PIN mem_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 256.950000 0.520000 257.050000 ;
    END
  END mem_in[98]
  PIN mem_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 254.950000 0.520000 255.050000 ;
    END
  END mem_in[97]
  PIN mem_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 252.950000 0.520000 253.050000 ;
    END
  END mem_in[96]
  PIN mem_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 250.950000 0.520000 251.050000 ;
    END
  END mem_in[95]
  PIN mem_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 248.950000 0.520000 249.050000 ;
    END
  END mem_in[94]
  PIN mem_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 246.950000 0.520000 247.050000 ;
    END
  END mem_in[93]
  PIN mem_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 244.950000 0.520000 245.050000 ;
    END
  END mem_in[92]
  PIN mem_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 242.950000 0.520000 243.050000 ;
    END
  END mem_in[91]
  PIN mem_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 240.950000 0.520000 241.050000 ;
    END
  END mem_in[90]
  PIN mem_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 238.950000 0.520000 239.050000 ;
    END
  END mem_in[89]
  PIN mem_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 236.950000 0.520000 237.050000 ;
    END
  END mem_in[88]
  PIN mem_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 234.950000 0.520000 235.050000 ;
    END
  END mem_in[87]
  PIN mem_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 232.950000 0.520000 233.050000 ;
    END
  END mem_in[86]
  PIN mem_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 230.950000 0.520000 231.050000 ;
    END
  END mem_in[85]
  PIN mem_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 228.950000 0.520000 229.050000 ;
    END
  END mem_in[84]
  PIN mem_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 226.950000 0.520000 227.050000 ;
    END
  END mem_in[83]
  PIN mem_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 224.950000 0.520000 225.050000 ;
    END
  END mem_in[82]
  PIN mem_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 222.950000 0.520000 223.050000 ;
    END
  END mem_in[81]
  PIN mem_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 220.950000 0.520000 221.050000 ;
    END
  END mem_in[80]
  PIN mem_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 218.950000 0.520000 219.050000 ;
    END
  END mem_in[79]
  PIN mem_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 216.950000 0.520000 217.050000 ;
    END
  END mem_in[78]
  PIN mem_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 214.950000 0.520000 215.050000 ;
    END
  END mem_in[77]
  PIN mem_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 212.950000 0.520000 213.050000 ;
    END
  END mem_in[76]
  PIN mem_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 210.950000 0.520000 211.050000 ;
    END
  END mem_in[75]
  PIN mem_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 208.950000 0.520000 209.050000 ;
    END
  END mem_in[74]
  PIN mem_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 206.950000 0.520000 207.050000 ;
    END
  END mem_in[73]
  PIN mem_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 204.950000 0.520000 205.050000 ;
    END
  END mem_in[72]
  PIN mem_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 202.950000 0.520000 203.050000 ;
    END
  END mem_in[71]
  PIN mem_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 200.950000 0.520000 201.050000 ;
    END
  END mem_in[70]
  PIN mem_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 198.950000 0.520000 199.050000 ;
    END
  END mem_in[69]
  PIN mem_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 196.950000 0.520000 197.050000 ;
    END
  END mem_in[68]
  PIN mem_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 194.950000 0.520000 195.050000 ;
    END
  END mem_in[67]
  PIN mem_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 192.950000 0.520000 193.050000 ;
    END
  END mem_in[66]
  PIN mem_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 190.950000 0.520000 191.050000 ;
    END
  END mem_in[65]
  PIN mem_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 188.950000 0.520000 189.050000 ;
    END
  END mem_in[64]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 186.950000 0.520000 187.050000 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 184.950000 0.520000 185.050000 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 182.950000 0.520000 183.050000 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 180.950000 0.520000 181.050000 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 178.950000 0.520000 179.050000 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 176.950000 0.520000 177.050000 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 174.950000 0.520000 175.050000 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 172.950000 0.520000 173.050000 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 170.950000 0.520000 171.050000 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 168.950000 0.520000 169.050000 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 166.950000 0.520000 167.050000 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 164.950000 0.520000 165.050000 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 162.950000 0.520000 163.050000 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 160.950000 0.520000 161.050000 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 158.950000 0.520000 159.050000 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 156.950000 0.520000 157.050000 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 154.950000 0.520000 155.050000 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 152.950000 0.520000 153.050000 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 150.950000 0.520000 151.050000 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 148.950000 0.520000 149.050000 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 146.950000 0.520000 147.050000 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 144.950000 0.520000 145.050000 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 142.950000 0.520000 143.050000 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 140.950000 0.520000 141.050000 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 138.950000 0.520000 139.050000 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 136.950000 0.520000 137.050000 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 134.950000 0.520000 135.050000 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 132.950000 0.520000 133.050000 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 130.950000 0.520000 131.050000 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 128.950000 0.520000 129.050000 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 126.950000 0.520000 127.050000 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 124.950000 0.520000 125.050000 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 122.950000 0.520000 123.050000 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 120.950000 0.520000 121.050000 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 118.950000 0.520000 119.050000 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 116.950000 0.520000 117.050000 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 114.950000 0.520000 115.050000 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 112.950000 0.520000 113.050000 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 110.950000 0.520000 111.050000 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 108.950000 0.520000 109.050000 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 106.950000 0.520000 107.050000 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 104.950000 0.520000 105.050000 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 102.950000 0.520000 103.050000 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 100.950000 0.520000 101.050000 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 98.950000 0.520000 99.050000 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 96.950000 0.520000 97.050000 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 94.950000 0.520000 95.050000 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 92.950000 0.520000 93.050000 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 90.950000 0.520000 91.050000 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 88.950000 0.520000 89.050000 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 86.950000 0.520000 87.050000 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 84.950000 0.520000 85.050000 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 82.950000 0.520000 83.050000 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 80.950000 0.520000 81.050000 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 78.950000 0.520000 79.050000 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 76.950000 0.520000 77.050000 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 74.950000 0.520000 75.050000 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 72.950000 0.520000 73.050000 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 70.950000 0.520000 71.050000 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 68.950000 0.520000 69.050000 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 66.950000 0.520000 67.050000 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 64.950000 0.520000 65.050000 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 62.950000 0.520000 63.050000 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 60.950000 0.520000 61.050000 ;
    END
  END mem_in[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 58.950000 0.520000 59.050000 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 56.950000 0.520000 57.050000 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 54.950000 0.520000 55.050000 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 52.950000 0.520000 53.050000 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 50.950000 0.520000 51.050000 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 48.950000 0.520000 49.050000 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 46.950000 0.520000 47.050000 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 44.950000 0.520000 45.050000 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 42.950000 0.520000 43.050000 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 40.950000 0.520000 41.050000 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 38.950000 0.520000 39.050000 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 36.950000 0.520000 37.050000 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 34.950000 0.520000 35.050000 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 32.950000 0.520000 33.050000 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 30.950000 0.520000 31.050000 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 28.950000 0.520000 29.050000 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 26.950000 0.520000 27.050000 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 316.950000 0.520000 317.050000 ;
    END
  END reset
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 350.050000 0.000000 350.150000 0.520000 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 352.050000 0.000000 352.150000 0.520000 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 354.050000 0.000000 354.150000 0.520000 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 356.050000 0.000000 356.150000 0.520000 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 358.050000 0.000000 358.150000 0.520000 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 360.050000 0.000000 360.150000 0.520000 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 362.050000 0.000000 362.150000 0.520000 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 364.050000 0.000000 364.150000 0.520000 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 366.050000 0.000000 366.150000 0.520000 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 368.050000 0.000000 368.150000 0.520000 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 370.050000 0.000000 370.150000 0.520000 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 372.050000 0.000000 372.150000 0.520000 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 374.050000 0.000000 374.150000 0.520000 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 376.050000 0.000000 376.150000 0.520000 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 378.050000 0.000000 378.150000 0.520000 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 380.050000 0.000000 380.150000 0.520000 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 382.050000 0.000000 382.150000 0.520000 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 384.050000 0.000000 384.150000 0.520000 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 386.050000 0.000000 386.150000 0.520000 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 388.050000 0.000000 388.150000 0.520000 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 390.050000 0.000000 390.150000 0.520000 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 392.050000 0.000000 392.150000 0.520000 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 394.050000 0.000000 394.150000 0.520000 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 396.050000 0.000000 396.150000 0.520000 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 398.050000 0.000000 398.150000 0.520000 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 400.050000 0.000000 400.150000 0.520000 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 402.050000 0.000000 402.150000 0.520000 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 404.050000 0.000000 404.150000 0.520000 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 406.050000 0.000000 406.150000 0.520000 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 408.050000 0.000000 408.150000 0.520000 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 410.050000 0.000000 410.150000 0.520000 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 412.050000 0.000000 412.150000 0.520000 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 414.050000 0.000000 414.150000 0.520000 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 416.050000 0.000000 416.150000 0.520000 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 418.050000 0.000000 418.150000 0.520000 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 420.050000 0.000000 420.150000 0.520000 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 422.050000 0.000000 422.150000 0.520000 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 424.050000 0.000000 424.150000 0.520000 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 426.050000 0.000000 426.150000 0.520000 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 428.050000 0.000000 428.150000 0.520000 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 430.050000 0.000000 430.150000 0.520000 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 432.050000 0.000000 432.150000 0.520000 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 434.050000 0.000000 434.150000 0.520000 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 436.050000 0.000000 436.150000 0.520000 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 438.050000 0.000000 438.150000 0.520000 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 440.050000 0.000000 440.150000 0.520000 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 442.050000 0.000000 442.150000 0.520000 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 444.050000 0.000000 444.150000 0.520000 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 446.050000 0.000000 446.150000 0.520000 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 448.050000 0.000000 448.150000 0.520000 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 450.050000 0.000000 450.150000 0.520000 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 452.050000 0.000000 452.150000 0.520000 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 454.050000 0.000000 454.150000 0.520000 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 456.050000 0.000000 456.150000 0.520000 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 458.050000 0.000000 458.150000 0.520000 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 460.050000 0.000000 460.150000 0.520000 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 462.050000 0.000000 462.150000 0.520000 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 464.050000 0.000000 464.150000 0.520000 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 466.050000 0.000000 466.150000 0.520000 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 468.050000 0.000000 468.150000 0.520000 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 470.050000 0.000000 470.150000 0.520000 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 472.050000 0.000000 472.150000 0.520000 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 474.050000 0.000000 474.150000 0.520000 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 476.050000 0.000000 476.150000 0.520000 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 478.050000 0.000000 478.150000 0.520000 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 480.050000 0.000000 480.150000 0.520000 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 482.050000 0.000000 482.150000 0.520000 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 484.050000 0.000000 484.150000 0.520000 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 486.050000 0.000000 486.150000 0.520000 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 488.050000 0.000000 488.150000 0.520000 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 490.050000 0.000000 490.150000 0.520000 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 492.050000 0.000000 492.150000 0.520000 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 494.050000 0.000000 494.150000 0.520000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 496.050000 0.000000 496.150000 0.520000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 498.050000 0.000000 498.150000 0.520000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 500.050000 0.000000 500.150000 0.520000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 502.050000 0.000000 502.150000 0.520000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 504.050000 0.000000 504.150000 0.520000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 506.050000 0.000000 506.150000 0.520000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 508.050000 0.000000 508.150000 0.520000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 510.050000 0.000000 510.150000 0.520000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 512.050000 0.000000 512.150000 0.520000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 514.050000 0.000000 514.150000 0.520000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 516.050000 0.000000 516.150000 0.520000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 518.050000 0.000000 518.150000 0.520000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 520.050000 0.000000 520.150000 0.520000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 522.050000 0.000000 522.150000 0.520000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 524.050000 0.000000 524.150000 0.520000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 526.050000 0.000000 526.150000 0.520000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 528.050000 0.000000 528.150000 0.520000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 530.050000 0.000000 530.150000 0.520000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 532.050000 0.000000 532.150000 0.520000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 534.050000 0.000000 534.150000 0.520000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 536.050000 0.000000 536.150000 0.520000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 538.050000 0.000000 538.150000 0.520000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 540.050000 0.000000 540.150000 0.520000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 542.050000 0.000000 542.150000 0.520000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 544.050000 0.000000 544.150000 0.520000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 546.050000 0.000000 546.150000 0.520000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 548.050000 0.000000 548.150000 0.520000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 550.050000 0.000000 550.150000 0.520000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 552.050000 0.000000 552.150000 0.520000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 554.050000 0.000000 554.150000 0.520000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 556.050000 0.000000 556.150000 0.520000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 558.050000 0.000000 558.150000 0.520000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 560.050000 0.000000 560.150000 0.520000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 562.050000 0.000000 562.150000 0.520000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 564.050000 0.000000 564.150000 0.520000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 566.050000 0.000000 566.150000 0.520000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 568.050000 0.000000 568.150000 0.520000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 570.050000 0.000000 570.150000 0.520000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 572.050000 0.000000 572.150000 0.520000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 574.050000 0.000000 574.150000 0.520000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 576.050000 0.000000 576.150000 0.520000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 578.050000 0.000000 578.150000 0.520000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 580.050000 0.000000 580.150000 0.520000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 582.050000 0.000000 582.150000 0.520000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 584.050000 0.000000 584.150000 0.520000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 586.050000 0.000000 586.150000 0.520000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 588.050000 0.000000 588.150000 0.520000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 590.050000 0.000000 590.150000 0.520000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 592.050000 0.000000 592.150000 0.520000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 594.050000 0.000000 594.150000 0.520000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 596.050000 0.000000 596.150000 0.520000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 598.050000 0.000000 598.150000 0.520000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 600.050000 0.000000 600.150000 0.520000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 602.050000 0.000000 602.150000 0.520000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 604.050000 0.000000 604.150000 0.520000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 606.050000 0.000000 606.150000 0.520000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 608.050000 0.000000 608.150000 0.520000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 610.050000 0.000000 610.150000 0.520000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 612.050000 0.000000 612.150000 0.520000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 614.050000 0.000000 614.150000 0.520000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 616.050000 0.000000 616.150000 0.520000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 618.050000 0.000000 618.150000 0.520000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 620.050000 0.000000 620.150000 0.520000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 622.050000 0.000000 622.150000 0.520000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 624.050000 0.000000 624.150000 0.520000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 626.050000 0.000000 626.150000 0.520000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 628.050000 0.000000 628.150000 0.520000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 630.050000 0.000000 630.150000 0.520000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 632.050000 0.000000 632.150000 0.520000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 634.050000 0.000000 634.150000 0.520000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 636.050000 0.000000 636.150000 0.520000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 638.050000 0.000000 638.150000 0.520000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 640.050000 0.000000 640.150000 0.520000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 642.050000 0.000000 642.150000 0.520000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 644.050000 0.000000 644.150000 0.520000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 646.050000 0.000000 646.150000 0.520000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 648.050000 0.000000 648.150000 0.520000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 650.050000 0.000000 650.150000 0.520000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 652.050000 0.000000 652.150000 0.520000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 654.050000 0.000000 654.150000 0.520000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 656.050000 0.000000 656.150000 0.520000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 658.050000 0.000000 658.150000 0.520000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 660.050000 0.000000 660.150000 0.520000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 662.050000 0.000000 662.150000 0.520000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 664.050000 0.000000 664.150000 0.520000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 666.050000 0.000000 666.150000 0.520000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 668.050000 0.000000 668.150000 0.520000 ;
    END
  END out[0]
  PIN sum_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 302.050000 0.000000 302.150000 0.520000 ;
    END
  END sum_out[23]
  PIN sum_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 304.050000 0.000000 304.150000 0.520000 ;
    END
  END sum_out[22]
  PIN sum_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 306.050000 0.000000 306.150000 0.520000 ;
    END
  END sum_out[21]
  PIN sum_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 308.050000 0.000000 308.150000 0.520000 ;
    END
  END sum_out[20]
  PIN sum_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 310.050000 0.000000 310.150000 0.520000 ;
    END
  END sum_out[19]
  PIN sum_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 312.050000 0.000000 312.150000 0.520000 ;
    END
  END sum_out[18]
  PIN sum_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 314.050000 0.000000 314.150000 0.520000 ;
    END
  END sum_out[17]
  PIN sum_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 316.050000 0.000000 316.150000 0.520000 ;
    END
  END sum_out[16]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 318.050000 0.000000 318.150000 0.520000 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 320.050000 0.000000 320.150000 0.520000 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 322.050000 0.000000 322.150000 0.520000 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 324.050000 0.000000 324.150000 0.520000 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 326.050000 0.000000 326.150000 0.520000 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 328.050000 0.000000 328.150000 0.520000 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 330.050000 0.000000 330.150000 0.520000 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.050000 0.000000 332.150000 0.520000 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 334.050000 0.000000 334.150000 0.520000 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 336.050000 0.000000 336.150000 0.520000 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 338.050000 0.000000 338.150000 0.520000 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 340.050000 0.000000 340.150000 0.520000 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 342.050000 0.000000 342.150000 0.520000 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 344.050000 0.000000 344.150000 0.520000 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 346.050000 0.000000 346.150000 0.520000 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 348.050000 0.000000 348.150000 0.520000 ;
    END
  END sum_out[0]
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 693.200000 689.600000 ;
    LAYER M2 ;
      RECT 0.000000 0.640000 693.200000 689.600000 ;
      RECT 668.250000 0.000000 693.200000 0.640000 ;
      RECT 666.250000 0.000000 667.950000 0.640000 ;
      RECT 664.250000 0.000000 665.950000 0.640000 ;
      RECT 662.250000 0.000000 663.950000 0.640000 ;
      RECT 660.250000 0.000000 661.950000 0.640000 ;
      RECT 658.250000 0.000000 659.950000 0.640000 ;
      RECT 656.250000 0.000000 657.950000 0.640000 ;
      RECT 654.250000 0.000000 655.950000 0.640000 ;
      RECT 652.250000 0.000000 653.950000 0.640000 ;
      RECT 650.250000 0.000000 651.950000 0.640000 ;
      RECT 648.250000 0.000000 649.950000 0.640000 ;
      RECT 646.250000 0.000000 647.950000 0.640000 ;
      RECT 644.250000 0.000000 645.950000 0.640000 ;
      RECT 642.250000 0.000000 643.950000 0.640000 ;
      RECT 640.250000 0.000000 641.950000 0.640000 ;
      RECT 638.250000 0.000000 639.950000 0.640000 ;
      RECT 636.250000 0.000000 637.950000 0.640000 ;
      RECT 634.250000 0.000000 635.950000 0.640000 ;
      RECT 632.250000 0.000000 633.950000 0.640000 ;
      RECT 630.250000 0.000000 631.950000 0.640000 ;
      RECT 628.250000 0.000000 629.950000 0.640000 ;
      RECT 626.250000 0.000000 627.950000 0.640000 ;
      RECT 624.250000 0.000000 625.950000 0.640000 ;
      RECT 622.250000 0.000000 623.950000 0.640000 ;
      RECT 620.250000 0.000000 621.950000 0.640000 ;
      RECT 618.250000 0.000000 619.950000 0.640000 ;
      RECT 616.250000 0.000000 617.950000 0.640000 ;
      RECT 614.250000 0.000000 615.950000 0.640000 ;
      RECT 612.250000 0.000000 613.950000 0.640000 ;
      RECT 610.250000 0.000000 611.950000 0.640000 ;
      RECT 608.250000 0.000000 609.950000 0.640000 ;
      RECT 606.250000 0.000000 607.950000 0.640000 ;
      RECT 604.250000 0.000000 605.950000 0.640000 ;
      RECT 602.250000 0.000000 603.950000 0.640000 ;
      RECT 600.250000 0.000000 601.950000 0.640000 ;
      RECT 598.250000 0.000000 599.950000 0.640000 ;
      RECT 596.250000 0.000000 597.950000 0.640000 ;
      RECT 594.250000 0.000000 595.950000 0.640000 ;
      RECT 592.250000 0.000000 593.950000 0.640000 ;
      RECT 590.250000 0.000000 591.950000 0.640000 ;
      RECT 588.250000 0.000000 589.950000 0.640000 ;
      RECT 586.250000 0.000000 587.950000 0.640000 ;
      RECT 584.250000 0.000000 585.950000 0.640000 ;
      RECT 582.250000 0.000000 583.950000 0.640000 ;
      RECT 580.250000 0.000000 581.950000 0.640000 ;
      RECT 578.250000 0.000000 579.950000 0.640000 ;
      RECT 576.250000 0.000000 577.950000 0.640000 ;
      RECT 574.250000 0.000000 575.950000 0.640000 ;
      RECT 572.250000 0.000000 573.950000 0.640000 ;
      RECT 570.250000 0.000000 571.950000 0.640000 ;
      RECT 568.250000 0.000000 569.950000 0.640000 ;
      RECT 566.250000 0.000000 567.950000 0.640000 ;
      RECT 564.250000 0.000000 565.950000 0.640000 ;
      RECT 562.250000 0.000000 563.950000 0.640000 ;
      RECT 560.250000 0.000000 561.950000 0.640000 ;
      RECT 558.250000 0.000000 559.950000 0.640000 ;
      RECT 556.250000 0.000000 557.950000 0.640000 ;
      RECT 554.250000 0.000000 555.950000 0.640000 ;
      RECT 552.250000 0.000000 553.950000 0.640000 ;
      RECT 550.250000 0.000000 551.950000 0.640000 ;
      RECT 548.250000 0.000000 549.950000 0.640000 ;
      RECT 546.250000 0.000000 547.950000 0.640000 ;
      RECT 544.250000 0.000000 545.950000 0.640000 ;
      RECT 542.250000 0.000000 543.950000 0.640000 ;
      RECT 540.250000 0.000000 541.950000 0.640000 ;
      RECT 538.250000 0.000000 539.950000 0.640000 ;
      RECT 536.250000 0.000000 537.950000 0.640000 ;
      RECT 534.250000 0.000000 535.950000 0.640000 ;
      RECT 532.250000 0.000000 533.950000 0.640000 ;
      RECT 530.250000 0.000000 531.950000 0.640000 ;
      RECT 528.250000 0.000000 529.950000 0.640000 ;
      RECT 526.250000 0.000000 527.950000 0.640000 ;
      RECT 524.250000 0.000000 525.950000 0.640000 ;
      RECT 522.250000 0.000000 523.950000 0.640000 ;
      RECT 520.250000 0.000000 521.950000 0.640000 ;
      RECT 518.250000 0.000000 519.950000 0.640000 ;
      RECT 516.250000 0.000000 517.950000 0.640000 ;
      RECT 514.250000 0.000000 515.950000 0.640000 ;
      RECT 512.250000 0.000000 513.950000 0.640000 ;
      RECT 510.250000 0.000000 511.950000 0.640000 ;
      RECT 508.250000 0.000000 509.950000 0.640000 ;
      RECT 506.250000 0.000000 507.950000 0.640000 ;
      RECT 504.250000 0.000000 505.950000 0.640000 ;
      RECT 502.250000 0.000000 503.950000 0.640000 ;
      RECT 500.250000 0.000000 501.950000 0.640000 ;
      RECT 498.250000 0.000000 499.950000 0.640000 ;
      RECT 496.250000 0.000000 497.950000 0.640000 ;
      RECT 494.250000 0.000000 495.950000 0.640000 ;
      RECT 492.250000 0.000000 493.950000 0.640000 ;
      RECT 490.250000 0.000000 491.950000 0.640000 ;
      RECT 488.250000 0.000000 489.950000 0.640000 ;
      RECT 486.250000 0.000000 487.950000 0.640000 ;
      RECT 484.250000 0.000000 485.950000 0.640000 ;
      RECT 482.250000 0.000000 483.950000 0.640000 ;
      RECT 480.250000 0.000000 481.950000 0.640000 ;
      RECT 478.250000 0.000000 479.950000 0.640000 ;
      RECT 476.250000 0.000000 477.950000 0.640000 ;
      RECT 474.250000 0.000000 475.950000 0.640000 ;
      RECT 472.250000 0.000000 473.950000 0.640000 ;
      RECT 470.250000 0.000000 471.950000 0.640000 ;
      RECT 468.250000 0.000000 469.950000 0.640000 ;
      RECT 466.250000 0.000000 467.950000 0.640000 ;
      RECT 464.250000 0.000000 465.950000 0.640000 ;
      RECT 462.250000 0.000000 463.950000 0.640000 ;
      RECT 460.250000 0.000000 461.950000 0.640000 ;
      RECT 458.250000 0.000000 459.950000 0.640000 ;
      RECT 456.250000 0.000000 457.950000 0.640000 ;
      RECT 454.250000 0.000000 455.950000 0.640000 ;
      RECT 452.250000 0.000000 453.950000 0.640000 ;
      RECT 450.250000 0.000000 451.950000 0.640000 ;
      RECT 448.250000 0.000000 449.950000 0.640000 ;
      RECT 446.250000 0.000000 447.950000 0.640000 ;
      RECT 444.250000 0.000000 445.950000 0.640000 ;
      RECT 442.250000 0.000000 443.950000 0.640000 ;
      RECT 440.250000 0.000000 441.950000 0.640000 ;
      RECT 438.250000 0.000000 439.950000 0.640000 ;
      RECT 436.250000 0.000000 437.950000 0.640000 ;
      RECT 434.250000 0.000000 435.950000 0.640000 ;
      RECT 432.250000 0.000000 433.950000 0.640000 ;
      RECT 430.250000 0.000000 431.950000 0.640000 ;
      RECT 428.250000 0.000000 429.950000 0.640000 ;
      RECT 426.250000 0.000000 427.950000 0.640000 ;
      RECT 424.250000 0.000000 425.950000 0.640000 ;
      RECT 422.250000 0.000000 423.950000 0.640000 ;
      RECT 420.250000 0.000000 421.950000 0.640000 ;
      RECT 418.250000 0.000000 419.950000 0.640000 ;
      RECT 416.250000 0.000000 417.950000 0.640000 ;
      RECT 414.250000 0.000000 415.950000 0.640000 ;
      RECT 412.250000 0.000000 413.950000 0.640000 ;
      RECT 410.250000 0.000000 411.950000 0.640000 ;
      RECT 408.250000 0.000000 409.950000 0.640000 ;
      RECT 406.250000 0.000000 407.950000 0.640000 ;
      RECT 404.250000 0.000000 405.950000 0.640000 ;
      RECT 402.250000 0.000000 403.950000 0.640000 ;
      RECT 400.250000 0.000000 401.950000 0.640000 ;
      RECT 398.250000 0.000000 399.950000 0.640000 ;
      RECT 396.250000 0.000000 397.950000 0.640000 ;
      RECT 394.250000 0.000000 395.950000 0.640000 ;
      RECT 392.250000 0.000000 393.950000 0.640000 ;
      RECT 390.250000 0.000000 391.950000 0.640000 ;
      RECT 388.250000 0.000000 389.950000 0.640000 ;
      RECT 386.250000 0.000000 387.950000 0.640000 ;
      RECT 384.250000 0.000000 385.950000 0.640000 ;
      RECT 382.250000 0.000000 383.950000 0.640000 ;
      RECT 380.250000 0.000000 381.950000 0.640000 ;
      RECT 378.250000 0.000000 379.950000 0.640000 ;
      RECT 376.250000 0.000000 377.950000 0.640000 ;
      RECT 374.250000 0.000000 375.950000 0.640000 ;
      RECT 372.250000 0.000000 373.950000 0.640000 ;
      RECT 370.250000 0.000000 371.950000 0.640000 ;
      RECT 368.250000 0.000000 369.950000 0.640000 ;
      RECT 366.250000 0.000000 367.950000 0.640000 ;
      RECT 364.250000 0.000000 365.950000 0.640000 ;
      RECT 362.250000 0.000000 363.950000 0.640000 ;
      RECT 360.250000 0.000000 361.950000 0.640000 ;
      RECT 358.250000 0.000000 359.950000 0.640000 ;
      RECT 356.250000 0.000000 357.950000 0.640000 ;
      RECT 354.250000 0.000000 355.950000 0.640000 ;
      RECT 352.250000 0.000000 353.950000 0.640000 ;
      RECT 350.250000 0.000000 351.950000 0.640000 ;
      RECT 348.250000 0.000000 349.950000 0.640000 ;
      RECT 346.250000 0.000000 347.950000 0.640000 ;
      RECT 344.250000 0.000000 345.950000 0.640000 ;
      RECT 342.250000 0.000000 343.950000 0.640000 ;
      RECT 340.250000 0.000000 341.950000 0.640000 ;
      RECT 338.250000 0.000000 339.950000 0.640000 ;
      RECT 336.250000 0.000000 337.950000 0.640000 ;
      RECT 334.250000 0.000000 335.950000 0.640000 ;
      RECT 332.250000 0.000000 333.950000 0.640000 ;
      RECT 330.250000 0.000000 331.950000 0.640000 ;
      RECT 328.250000 0.000000 329.950000 0.640000 ;
      RECT 326.250000 0.000000 327.950000 0.640000 ;
      RECT 324.250000 0.000000 325.950000 0.640000 ;
      RECT 322.250000 0.000000 323.950000 0.640000 ;
      RECT 320.250000 0.000000 321.950000 0.640000 ;
      RECT 318.250000 0.000000 319.950000 0.640000 ;
      RECT 316.250000 0.000000 317.950000 0.640000 ;
      RECT 314.250000 0.000000 315.950000 0.640000 ;
      RECT 312.250000 0.000000 313.950000 0.640000 ;
      RECT 310.250000 0.000000 311.950000 0.640000 ;
      RECT 308.250000 0.000000 309.950000 0.640000 ;
      RECT 306.250000 0.000000 307.950000 0.640000 ;
      RECT 304.250000 0.000000 305.950000 0.640000 ;
      RECT 302.250000 0.000000 303.950000 0.640000 ;
      RECT 0.000000 0.000000 301.950000 0.640000 ;
    LAYER M3 ;
      RECT 0.000000 317.150000 693.200000 689.600000 ;
      RECT 0.640000 316.850000 693.200000 317.150000 ;
      RECT 0.000000 315.150000 693.200000 316.850000 ;
      RECT 0.640000 314.850000 693.200000 315.150000 ;
      RECT 0.000000 313.150000 693.200000 314.850000 ;
      RECT 0.640000 312.850000 693.200000 313.150000 ;
      RECT 0.000000 311.150000 693.200000 312.850000 ;
      RECT 0.640000 310.850000 693.200000 311.150000 ;
      RECT 0.000000 309.150000 693.200000 310.850000 ;
      RECT 0.640000 308.850000 693.200000 309.150000 ;
      RECT 0.000000 307.150000 693.200000 308.850000 ;
      RECT 0.640000 306.850000 693.200000 307.150000 ;
      RECT 0.000000 305.150000 693.200000 306.850000 ;
      RECT 0.640000 304.850000 693.200000 305.150000 ;
      RECT 0.000000 303.150000 693.200000 304.850000 ;
      RECT 0.640000 302.850000 693.200000 303.150000 ;
      RECT 0.000000 301.150000 693.200000 302.850000 ;
      RECT 0.640000 300.850000 693.200000 301.150000 ;
      RECT 0.000000 299.150000 693.200000 300.850000 ;
      RECT 0.640000 298.850000 693.200000 299.150000 ;
      RECT 0.000000 297.150000 693.200000 298.850000 ;
      RECT 0.640000 296.850000 693.200000 297.150000 ;
      RECT 0.000000 295.150000 693.200000 296.850000 ;
      RECT 0.640000 294.850000 693.200000 295.150000 ;
      RECT 0.000000 293.150000 693.200000 294.850000 ;
      RECT 0.640000 292.850000 693.200000 293.150000 ;
      RECT 0.000000 291.150000 693.200000 292.850000 ;
      RECT 0.640000 290.850000 693.200000 291.150000 ;
      RECT 0.000000 289.150000 693.200000 290.850000 ;
      RECT 0.640000 288.850000 693.200000 289.150000 ;
      RECT 0.000000 287.150000 693.200000 288.850000 ;
      RECT 0.640000 286.850000 693.200000 287.150000 ;
      RECT 0.000000 285.150000 693.200000 286.850000 ;
      RECT 0.640000 284.850000 693.200000 285.150000 ;
      RECT 0.000000 283.150000 693.200000 284.850000 ;
      RECT 0.640000 282.850000 693.200000 283.150000 ;
      RECT 0.000000 281.150000 693.200000 282.850000 ;
      RECT 0.640000 280.850000 693.200000 281.150000 ;
      RECT 0.000000 279.150000 693.200000 280.850000 ;
      RECT 0.640000 278.850000 693.200000 279.150000 ;
      RECT 0.000000 277.150000 693.200000 278.850000 ;
      RECT 0.640000 276.850000 693.200000 277.150000 ;
      RECT 0.000000 275.150000 693.200000 276.850000 ;
      RECT 0.640000 274.850000 693.200000 275.150000 ;
      RECT 0.000000 273.150000 693.200000 274.850000 ;
      RECT 0.640000 272.850000 693.200000 273.150000 ;
      RECT 0.000000 271.150000 693.200000 272.850000 ;
      RECT 0.640000 270.850000 693.200000 271.150000 ;
      RECT 0.000000 269.150000 693.200000 270.850000 ;
      RECT 0.640000 268.850000 693.200000 269.150000 ;
      RECT 0.000000 267.150000 693.200000 268.850000 ;
      RECT 0.640000 266.850000 693.200000 267.150000 ;
      RECT 0.000000 265.150000 693.200000 266.850000 ;
      RECT 0.640000 264.850000 693.200000 265.150000 ;
      RECT 0.000000 263.150000 693.200000 264.850000 ;
      RECT 0.640000 262.850000 693.200000 263.150000 ;
      RECT 0.000000 261.150000 693.200000 262.850000 ;
      RECT 0.640000 260.850000 693.200000 261.150000 ;
      RECT 0.000000 259.150000 693.200000 260.850000 ;
      RECT 0.640000 258.850000 693.200000 259.150000 ;
      RECT 0.000000 257.150000 693.200000 258.850000 ;
      RECT 0.640000 256.850000 693.200000 257.150000 ;
      RECT 0.000000 255.150000 693.200000 256.850000 ;
      RECT 0.640000 254.850000 693.200000 255.150000 ;
      RECT 0.000000 253.150000 693.200000 254.850000 ;
      RECT 0.640000 252.850000 693.200000 253.150000 ;
      RECT 0.000000 251.150000 693.200000 252.850000 ;
      RECT 0.640000 250.850000 693.200000 251.150000 ;
      RECT 0.000000 249.150000 693.200000 250.850000 ;
      RECT 0.640000 248.850000 693.200000 249.150000 ;
      RECT 0.000000 247.150000 693.200000 248.850000 ;
      RECT 0.640000 246.850000 693.200000 247.150000 ;
      RECT 0.000000 245.150000 693.200000 246.850000 ;
      RECT 0.640000 244.850000 693.200000 245.150000 ;
      RECT 0.000000 243.150000 693.200000 244.850000 ;
      RECT 0.640000 242.850000 693.200000 243.150000 ;
      RECT 0.000000 241.150000 693.200000 242.850000 ;
      RECT 0.640000 240.850000 693.200000 241.150000 ;
      RECT 0.000000 239.150000 693.200000 240.850000 ;
      RECT 0.640000 238.850000 693.200000 239.150000 ;
      RECT 0.000000 237.150000 693.200000 238.850000 ;
      RECT 0.640000 236.850000 693.200000 237.150000 ;
      RECT 0.000000 235.150000 693.200000 236.850000 ;
      RECT 0.640000 234.850000 693.200000 235.150000 ;
      RECT 0.000000 233.150000 693.200000 234.850000 ;
      RECT 0.640000 232.850000 693.200000 233.150000 ;
      RECT 0.000000 231.150000 693.200000 232.850000 ;
      RECT 0.640000 230.850000 693.200000 231.150000 ;
      RECT 0.000000 229.150000 693.200000 230.850000 ;
      RECT 0.640000 228.850000 693.200000 229.150000 ;
      RECT 0.000000 227.150000 693.200000 228.850000 ;
      RECT 0.640000 226.850000 693.200000 227.150000 ;
      RECT 0.000000 225.150000 693.200000 226.850000 ;
      RECT 0.640000 224.850000 693.200000 225.150000 ;
      RECT 0.000000 223.150000 693.200000 224.850000 ;
      RECT 0.640000 222.850000 693.200000 223.150000 ;
      RECT 0.000000 221.150000 693.200000 222.850000 ;
      RECT 0.640000 220.850000 693.200000 221.150000 ;
      RECT 0.000000 219.150000 693.200000 220.850000 ;
      RECT 0.640000 218.850000 693.200000 219.150000 ;
      RECT 0.000000 217.150000 693.200000 218.850000 ;
      RECT 0.640000 216.850000 693.200000 217.150000 ;
      RECT 0.000000 215.150000 693.200000 216.850000 ;
      RECT 0.640000 214.850000 693.200000 215.150000 ;
      RECT 0.000000 213.150000 693.200000 214.850000 ;
      RECT 0.640000 212.850000 693.200000 213.150000 ;
      RECT 0.000000 211.150000 693.200000 212.850000 ;
      RECT 0.640000 210.850000 693.200000 211.150000 ;
      RECT 0.000000 209.150000 693.200000 210.850000 ;
      RECT 0.640000 208.850000 693.200000 209.150000 ;
      RECT 0.000000 207.150000 693.200000 208.850000 ;
      RECT 0.640000 206.850000 693.200000 207.150000 ;
      RECT 0.000000 205.150000 693.200000 206.850000 ;
      RECT 0.640000 204.850000 693.200000 205.150000 ;
      RECT 0.000000 203.150000 693.200000 204.850000 ;
      RECT 0.640000 202.850000 693.200000 203.150000 ;
      RECT 0.000000 201.150000 693.200000 202.850000 ;
      RECT 0.640000 200.850000 693.200000 201.150000 ;
      RECT 0.000000 199.150000 693.200000 200.850000 ;
      RECT 0.640000 198.850000 693.200000 199.150000 ;
      RECT 0.000000 197.150000 693.200000 198.850000 ;
      RECT 0.640000 196.850000 693.200000 197.150000 ;
      RECT 0.000000 195.150000 693.200000 196.850000 ;
      RECT 0.640000 194.850000 693.200000 195.150000 ;
      RECT 0.000000 193.150000 693.200000 194.850000 ;
      RECT 0.640000 192.850000 693.200000 193.150000 ;
      RECT 0.000000 191.150000 693.200000 192.850000 ;
      RECT 0.640000 190.850000 693.200000 191.150000 ;
      RECT 0.000000 189.150000 693.200000 190.850000 ;
      RECT 0.640000 188.850000 693.200000 189.150000 ;
      RECT 0.000000 187.150000 693.200000 188.850000 ;
      RECT 0.640000 186.850000 693.200000 187.150000 ;
      RECT 0.000000 185.150000 693.200000 186.850000 ;
      RECT 0.640000 184.850000 693.200000 185.150000 ;
      RECT 0.000000 183.150000 693.200000 184.850000 ;
      RECT 0.640000 182.850000 693.200000 183.150000 ;
      RECT 0.000000 181.150000 693.200000 182.850000 ;
      RECT 0.640000 180.850000 693.200000 181.150000 ;
      RECT 0.000000 179.150000 693.200000 180.850000 ;
      RECT 0.640000 178.850000 693.200000 179.150000 ;
      RECT 0.000000 177.150000 693.200000 178.850000 ;
      RECT 0.640000 176.850000 693.200000 177.150000 ;
      RECT 0.000000 175.150000 693.200000 176.850000 ;
      RECT 0.640000 174.850000 693.200000 175.150000 ;
      RECT 0.000000 173.150000 693.200000 174.850000 ;
      RECT 0.640000 172.850000 693.200000 173.150000 ;
      RECT 0.000000 171.150000 693.200000 172.850000 ;
      RECT 0.640000 170.850000 693.200000 171.150000 ;
      RECT 0.000000 169.150000 693.200000 170.850000 ;
      RECT 0.640000 168.850000 693.200000 169.150000 ;
      RECT 0.000000 167.150000 693.200000 168.850000 ;
      RECT 0.640000 166.850000 693.200000 167.150000 ;
      RECT 0.000000 165.150000 693.200000 166.850000 ;
      RECT 0.640000 164.850000 693.200000 165.150000 ;
      RECT 0.000000 163.150000 693.200000 164.850000 ;
      RECT 0.640000 162.850000 693.200000 163.150000 ;
      RECT 0.000000 161.150000 693.200000 162.850000 ;
      RECT 0.640000 160.850000 693.200000 161.150000 ;
      RECT 0.000000 159.150000 693.200000 160.850000 ;
      RECT 0.640000 158.850000 693.200000 159.150000 ;
      RECT 0.000000 157.150000 693.200000 158.850000 ;
      RECT 0.640000 156.850000 693.200000 157.150000 ;
      RECT 0.000000 155.150000 693.200000 156.850000 ;
      RECT 0.640000 154.850000 693.200000 155.150000 ;
      RECT 0.000000 153.150000 693.200000 154.850000 ;
      RECT 0.640000 152.850000 693.200000 153.150000 ;
      RECT 0.000000 151.150000 693.200000 152.850000 ;
      RECT 0.640000 150.850000 693.200000 151.150000 ;
      RECT 0.000000 149.150000 693.200000 150.850000 ;
      RECT 0.640000 148.850000 693.200000 149.150000 ;
      RECT 0.000000 147.150000 693.200000 148.850000 ;
      RECT 0.640000 146.850000 693.200000 147.150000 ;
      RECT 0.000000 145.150000 693.200000 146.850000 ;
      RECT 0.640000 144.850000 693.200000 145.150000 ;
      RECT 0.000000 143.150000 693.200000 144.850000 ;
      RECT 0.640000 142.850000 693.200000 143.150000 ;
      RECT 0.000000 141.150000 693.200000 142.850000 ;
      RECT 0.640000 140.850000 693.200000 141.150000 ;
      RECT 0.000000 139.150000 693.200000 140.850000 ;
      RECT 0.640000 138.850000 693.200000 139.150000 ;
      RECT 0.000000 137.150000 693.200000 138.850000 ;
      RECT 0.640000 136.850000 693.200000 137.150000 ;
      RECT 0.000000 135.150000 693.200000 136.850000 ;
      RECT 0.640000 134.850000 693.200000 135.150000 ;
      RECT 0.000000 133.150000 693.200000 134.850000 ;
      RECT 0.640000 132.850000 693.200000 133.150000 ;
      RECT 0.000000 131.150000 693.200000 132.850000 ;
      RECT 0.640000 130.850000 693.200000 131.150000 ;
      RECT 0.000000 129.150000 693.200000 130.850000 ;
      RECT 0.640000 128.850000 693.200000 129.150000 ;
      RECT 0.000000 127.150000 693.200000 128.850000 ;
      RECT 0.640000 126.850000 693.200000 127.150000 ;
      RECT 0.000000 125.150000 693.200000 126.850000 ;
      RECT 0.640000 124.850000 693.200000 125.150000 ;
      RECT 0.000000 123.150000 693.200000 124.850000 ;
      RECT 0.640000 122.850000 693.200000 123.150000 ;
      RECT 0.000000 121.150000 693.200000 122.850000 ;
      RECT 0.640000 120.850000 693.200000 121.150000 ;
      RECT 0.000000 119.150000 693.200000 120.850000 ;
      RECT 0.640000 118.850000 693.200000 119.150000 ;
      RECT 0.000000 117.150000 693.200000 118.850000 ;
      RECT 0.640000 116.850000 693.200000 117.150000 ;
      RECT 0.000000 115.150000 693.200000 116.850000 ;
      RECT 0.640000 114.850000 693.200000 115.150000 ;
      RECT 0.000000 113.150000 693.200000 114.850000 ;
      RECT 0.640000 112.850000 693.200000 113.150000 ;
      RECT 0.000000 111.150000 693.200000 112.850000 ;
      RECT 0.640000 110.850000 693.200000 111.150000 ;
      RECT 0.000000 109.150000 693.200000 110.850000 ;
      RECT 0.640000 108.850000 693.200000 109.150000 ;
      RECT 0.000000 107.150000 693.200000 108.850000 ;
      RECT 0.640000 106.850000 693.200000 107.150000 ;
      RECT 0.000000 105.150000 693.200000 106.850000 ;
      RECT 0.640000 104.850000 693.200000 105.150000 ;
      RECT 0.000000 103.150000 693.200000 104.850000 ;
      RECT 0.640000 102.850000 693.200000 103.150000 ;
      RECT 0.000000 101.150000 693.200000 102.850000 ;
      RECT 0.640000 100.850000 693.200000 101.150000 ;
      RECT 0.000000 99.150000 693.200000 100.850000 ;
      RECT 0.640000 98.850000 693.200000 99.150000 ;
      RECT 0.000000 97.150000 693.200000 98.850000 ;
      RECT 0.640000 96.850000 693.200000 97.150000 ;
      RECT 0.000000 95.150000 693.200000 96.850000 ;
      RECT 0.640000 94.850000 693.200000 95.150000 ;
      RECT 0.000000 93.150000 693.200000 94.850000 ;
      RECT 0.640000 92.850000 693.200000 93.150000 ;
      RECT 0.000000 91.150000 693.200000 92.850000 ;
      RECT 0.640000 90.850000 693.200000 91.150000 ;
      RECT 0.000000 89.150000 693.200000 90.850000 ;
      RECT 0.640000 88.850000 693.200000 89.150000 ;
      RECT 0.000000 87.150000 693.200000 88.850000 ;
      RECT 0.640000 86.850000 693.200000 87.150000 ;
      RECT 0.000000 85.150000 693.200000 86.850000 ;
      RECT 0.640000 84.850000 693.200000 85.150000 ;
      RECT 0.000000 83.150000 693.200000 84.850000 ;
      RECT 0.640000 82.850000 693.200000 83.150000 ;
      RECT 0.000000 81.150000 693.200000 82.850000 ;
      RECT 0.640000 80.850000 693.200000 81.150000 ;
      RECT 0.000000 79.150000 693.200000 80.850000 ;
      RECT 0.640000 78.850000 693.200000 79.150000 ;
      RECT 0.000000 77.150000 693.200000 78.850000 ;
      RECT 0.640000 76.850000 693.200000 77.150000 ;
      RECT 0.000000 75.150000 693.200000 76.850000 ;
      RECT 0.640000 74.850000 693.200000 75.150000 ;
      RECT 0.000000 73.150000 693.200000 74.850000 ;
      RECT 0.640000 72.850000 693.200000 73.150000 ;
      RECT 0.000000 71.150000 693.200000 72.850000 ;
      RECT 0.640000 70.850000 693.200000 71.150000 ;
      RECT 0.000000 69.150000 693.200000 70.850000 ;
      RECT 0.640000 68.850000 693.200000 69.150000 ;
      RECT 0.000000 67.150000 693.200000 68.850000 ;
      RECT 0.640000 66.850000 693.200000 67.150000 ;
      RECT 0.000000 65.150000 693.200000 66.850000 ;
      RECT 0.640000 64.850000 693.200000 65.150000 ;
      RECT 0.000000 63.150000 693.200000 64.850000 ;
      RECT 0.640000 62.850000 693.200000 63.150000 ;
      RECT 0.000000 61.150000 693.200000 62.850000 ;
      RECT 0.640000 60.850000 693.200000 61.150000 ;
      RECT 0.000000 59.150000 693.200000 60.850000 ;
      RECT 0.640000 58.850000 693.200000 59.150000 ;
      RECT 0.000000 57.150000 693.200000 58.850000 ;
      RECT 0.640000 56.850000 693.200000 57.150000 ;
      RECT 0.000000 55.150000 693.200000 56.850000 ;
      RECT 0.640000 54.850000 693.200000 55.150000 ;
      RECT 0.000000 53.150000 693.200000 54.850000 ;
      RECT 0.640000 52.850000 693.200000 53.150000 ;
      RECT 0.000000 51.150000 693.200000 52.850000 ;
      RECT 0.640000 50.850000 693.200000 51.150000 ;
      RECT 0.000000 49.150000 693.200000 50.850000 ;
      RECT 0.640000 48.850000 693.200000 49.150000 ;
      RECT 0.000000 47.150000 693.200000 48.850000 ;
      RECT 0.640000 46.850000 693.200000 47.150000 ;
      RECT 0.000000 45.150000 693.200000 46.850000 ;
      RECT 0.640000 44.850000 693.200000 45.150000 ;
      RECT 0.000000 43.150000 693.200000 44.850000 ;
      RECT 0.640000 42.850000 693.200000 43.150000 ;
      RECT 0.000000 41.150000 693.200000 42.850000 ;
      RECT 0.640000 40.850000 693.200000 41.150000 ;
      RECT 0.000000 39.150000 693.200000 40.850000 ;
      RECT 0.640000 38.850000 693.200000 39.150000 ;
      RECT 0.000000 37.150000 693.200000 38.850000 ;
      RECT 0.640000 36.850000 693.200000 37.150000 ;
      RECT 0.000000 35.150000 693.200000 36.850000 ;
      RECT 0.640000 34.850000 693.200000 35.150000 ;
      RECT 0.000000 33.150000 693.200000 34.850000 ;
      RECT 0.640000 32.850000 693.200000 33.150000 ;
      RECT 0.000000 31.150000 693.200000 32.850000 ;
      RECT 0.640000 30.850000 693.200000 31.150000 ;
      RECT 0.000000 29.150000 693.200000 30.850000 ;
      RECT 0.640000 28.850000 693.200000 29.150000 ;
      RECT 0.000000 27.150000 693.200000 28.850000 ;
      RECT 0.640000 26.850000 693.200000 27.150000 ;
      RECT 0.000000 25.150000 693.200000 26.850000 ;
      RECT 0.640000 24.850000 693.200000 25.150000 ;
      RECT 0.000000 0.000000 693.200000 24.850000 ;
    LAYER M4 ;
      RECT 0.000000 0.000000 693.200000 689.600000 ;
    LAYER M5 ;
      RECT 0.000000 0.000000 693.200000 689.600000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 693.200000 689.600000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 693.200000 689.600000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 693.200000 689.600000 ;
  END
END fullchip

END LIBRARY
