##
## LEF for PtnCells ;
## created by Innovus v19.17-s077_1 on Sun Mar 19 21:12:51 2023
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fullchip
  CLASS BLOCK ;
  SIZE 473.800000 BY 473.600000 ;
  FOREIGN fullchip 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 9.950000 0.520000 10.050000 ;
    END
  END clk
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 414.950000 0.520000 415.050000 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 409.950000 0.520000 410.050000 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 404.950000 0.520000 405.050000 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 399.950000 0.520000 400.050000 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 394.950000 0.520000 395.050000 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 389.950000 0.520000 390.050000 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 384.950000 0.520000 385.050000 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 379.950000 0.520000 380.050000 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 374.950000 0.520000 375.050000 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 369.950000 0.520000 370.050000 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 364.950000 0.520000 365.050000 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 359.950000 0.520000 360.050000 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 354.950000 0.520000 355.050000 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 349.950000 0.520000 350.050000 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 344.950000 0.520000 345.050000 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 339.950000 0.520000 340.050000 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 334.950000 0.520000 335.050000 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 329.950000 0.520000 330.050000 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 324.950000 0.520000 325.050000 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 319.950000 0.520000 320.050000 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 314.950000 0.520000 315.050000 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 309.950000 0.520000 310.050000 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 304.950000 0.520000 305.050000 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 299.950000 0.520000 300.050000 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 294.950000 0.520000 295.050000 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 289.950000 0.520000 290.050000 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 284.950000 0.520000 285.050000 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 279.950000 0.520000 280.050000 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 274.950000 0.520000 275.050000 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 269.950000 0.520000 270.050000 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 264.950000 0.520000 265.050000 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 259.950000 0.520000 260.050000 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 254.950000 0.520000 255.050000 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 249.950000 0.520000 250.050000 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 244.950000 0.520000 245.050000 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 239.950000 0.520000 240.050000 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 234.950000 0.520000 235.050000 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 229.950000 0.520000 230.050000 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 224.950000 0.520000 225.050000 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 219.950000 0.520000 220.050000 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 214.950000 0.520000 215.050000 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 209.950000 0.520000 210.050000 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 204.950000 0.520000 205.050000 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 199.950000 0.520000 200.050000 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 194.950000 0.520000 195.050000 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 189.950000 0.520000 190.050000 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 184.950000 0.520000 185.050000 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 179.950000 0.520000 180.050000 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 174.950000 0.520000 175.050000 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 169.950000 0.520000 170.050000 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 164.950000 0.520000 165.050000 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 159.950000 0.520000 160.050000 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 154.950000 0.520000 155.050000 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 149.950000 0.520000 150.050000 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 144.950000 0.520000 145.050000 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 139.950000 0.520000 140.050000 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 134.950000 0.520000 135.050000 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 129.950000 0.520000 130.050000 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 124.950000 0.520000 125.050000 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 119.950000 0.520000 120.050000 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 114.950000 0.520000 115.050000 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 109.950000 0.520000 110.050000 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 104.950000 0.520000 105.050000 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 99.950000 0.520000 100.050000 ;
    END
  END mem_in[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 94.950000 0.520000 95.050000 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 89.950000 0.520000 90.050000 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 84.950000 0.520000 85.050000 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 79.950000 0.520000 80.050000 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 74.950000 0.520000 75.050000 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 69.950000 0.520000 70.050000 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 64.950000 0.520000 65.050000 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 59.950000 0.520000 60.050000 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 54.950000 0.520000 55.050000 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 49.950000 0.520000 50.050000 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 44.950000 0.520000 45.050000 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 39.950000 0.520000 40.050000 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 34.950000 0.520000 35.050000 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 29.950000 0.520000 30.050000 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 24.950000 0.520000 25.050000 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 19.950000 0.520000 20.050000 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 14.950000 0.520000 15.050000 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 419.950000 0.520000 420.050000 ;
    END
  END reset
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.650000 0.000000 178.750000 0.520000 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 181.650000 0.000000 181.750000 0.520000 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 184.650000 0.000000 184.750000 0.520000 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 187.650000 0.000000 187.750000 0.520000 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.650000 0.000000 190.750000 0.520000 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 193.650000 0.000000 193.750000 0.520000 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.650000 0.000000 196.750000 0.520000 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 199.650000 0.000000 199.750000 0.520000 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 202.650000 0.000000 202.750000 0.520000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.650000 0.000000 205.750000 0.520000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 208.650000 0.000000 208.750000 0.520000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.650000 0.000000 211.750000 0.520000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 214.650000 0.000000 214.750000 0.520000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 217.650000 0.000000 217.750000 0.520000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 220.650000 0.000000 220.750000 0.520000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 223.650000 0.000000 223.750000 0.520000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.650000 0.000000 226.750000 0.520000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 229.650000 0.000000 229.750000 0.520000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 232.650000 0.000000 232.750000 0.520000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 235.650000 0.000000 235.750000 0.520000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 238.650000 0.000000 238.750000 0.520000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 241.650000 0.000000 241.750000 0.520000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 244.650000 0.000000 244.750000 0.520000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 247.650000 0.000000 247.750000 0.520000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 250.650000 0.000000 250.750000 0.520000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 253.650000 0.000000 253.750000 0.520000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 256.650000 0.000000 256.750000 0.520000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 259.650000 0.000000 259.750000 0.520000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 262.650000 0.000000 262.750000 0.520000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 265.650000 0.000000 265.750000 0.520000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 268.650000 0.000000 268.750000 0.520000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 271.650000 0.000000 271.750000 0.520000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 274.650000 0.000000 274.750000 0.520000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 277.650000 0.000000 277.750000 0.520000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 280.650000 0.000000 280.750000 0.520000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 283.650000 0.000000 283.750000 0.520000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 286.650000 0.000000 286.750000 0.520000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 289.650000 0.000000 289.750000 0.520000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 292.650000 0.000000 292.750000 0.520000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 295.650000 0.000000 295.750000 0.520000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 298.650000 0.000000 298.750000 0.520000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 301.650000 0.000000 301.750000 0.520000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 304.650000 0.000000 304.750000 0.520000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 307.650000 0.000000 307.750000 0.520000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 310.650000 0.000000 310.750000 0.520000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 313.650000 0.000000 313.750000 0.520000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 316.650000 0.000000 316.750000 0.520000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 319.650000 0.000000 319.750000 0.520000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 322.650000 0.000000 322.750000 0.520000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 325.650000 0.000000 325.750000 0.520000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 328.650000 0.000000 328.750000 0.520000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 331.650000 0.000000 331.750000 0.520000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 334.650000 0.000000 334.750000 0.520000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 337.650000 0.000000 337.750000 0.520000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 340.650000 0.000000 340.750000 0.520000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 343.650000 0.000000 343.750000 0.520000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 346.650000 0.000000 346.750000 0.520000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 349.650000 0.000000 349.750000 0.520000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 352.650000 0.000000 352.750000 0.520000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 355.650000 0.000000 355.750000 0.520000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 358.650000 0.000000 358.750000 0.520000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 361.650000 0.000000 361.750000 0.520000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 364.650000 0.000000 364.750000 0.520000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 367.650000 0.000000 367.750000 0.520000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 370.650000 0.000000 370.750000 0.520000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 373.650000 0.000000 373.750000 0.520000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 376.650000 0.000000 376.750000 0.520000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 379.650000 0.000000 379.750000 0.520000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 382.650000 0.000000 382.750000 0.520000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 385.650000 0.000000 385.750000 0.520000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 388.650000 0.000000 388.750000 0.520000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 391.650000 0.000000 391.750000 0.520000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 394.650000 0.000000 394.750000 0.520000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 397.650000 0.000000 397.750000 0.520000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 400.650000 0.000000 400.750000 0.520000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 403.650000 0.000000 403.750000 0.520000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 406.650000 0.000000 406.750000 0.520000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 409.650000 0.000000 409.750000 0.520000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 412.650000 0.000000 412.750000 0.520000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 415.650000 0.000000 415.750000 0.520000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 418.650000 0.000000 418.750000 0.520000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 421.650000 0.000000 421.750000 0.520000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 424.650000 0.000000 424.750000 0.520000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 427.650000 0.000000 427.750000 0.520000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 430.650000 0.000000 430.750000 0.520000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 433.650000 0.000000 433.750000 0.520000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 436.650000 0.000000 436.750000 0.520000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 439.650000 0.000000 439.750000 0.520000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 442.650000 0.000000 442.750000 0.520000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 445.650000 0.000000 445.750000 0.520000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 448.650000 0.000000 448.750000 0.520000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 451.650000 0.000000 451.750000 0.520000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 454.650000 0.000000 454.750000 0.520000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 457.650000 0.000000 457.750000 0.520000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 460.650000 0.000000 460.750000 0.520000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 463.650000 0.000000 463.750000 0.520000 ;
    END
  END out[0]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.650000 0.000000 130.750000 0.520000 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.650000 0.000000 133.750000 0.520000 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.650000 0.000000 136.750000 0.520000 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.650000 0.000000 139.750000 0.520000 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.650000 0.000000 142.750000 0.520000 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.650000 0.000000 145.750000 0.520000 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.650000 0.000000 148.750000 0.520000 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 151.650000 0.000000 151.750000 0.520000 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.650000 0.000000 154.750000 0.520000 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.650000 0.000000 157.750000 0.520000 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.650000 0.000000 160.750000 0.520000 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 163.650000 0.000000 163.750000 0.520000 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 166.650000 0.000000 166.750000 0.520000 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 169.650000 0.000000 169.750000 0.520000 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 172.650000 0.000000 172.750000 0.520000 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.650000 0.000000 175.750000 0.520000 ;
    END
  END sum_out[0]
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 473.800000 473.600000 ;
    LAYER M2 ;
      RECT 0.000000 0.640000 473.800000 473.600000 ;
      RECT 463.850000 0.000000 473.800000 0.640000 ;
      RECT 460.850000 0.000000 463.550000 0.640000 ;
      RECT 457.850000 0.000000 460.550000 0.640000 ;
      RECT 454.850000 0.000000 457.550000 0.640000 ;
      RECT 451.850000 0.000000 454.550000 0.640000 ;
      RECT 448.850000 0.000000 451.550000 0.640000 ;
      RECT 445.850000 0.000000 448.550000 0.640000 ;
      RECT 442.850000 0.000000 445.550000 0.640000 ;
      RECT 439.850000 0.000000 442.550000 0.640000 ;
      RECT 436.850000 0.000000 439.550000 0.640000 ;
      RECT 433.850000 0.000000 436.550000 0.640000 ;
      RECT 430.850000 0.000000 433.550000 0.640000 ;
      RECT 427.850000 0.000000 430.550000 0.640000 ;
      RECT 424.850000 0.000000 427.550000 0.640000 ;
      RECT 421.850000 0.000000 424.550000 0.640000 ;
      RECT 418.850000 0.000000 421.550000 0.640000 ;
      RECT 415.850000 0.000000 418.550000 0.640000 ;
      RECT 412.850000 0.000000 415.550000 0.640000 ;
      RECT 409.850000 0.000000 412.550000 0.640000 ;
      RECT 406.850000 0.000000 409.550000 0.640000 ;
      RECT 403.850000 0.000000 406.550000 0.640000 ;
      RECT 400.850000 0.000000 403.550000 0.640000 ;
      RECT 397.850000 0.000000 400.550000 0.640000 ;
      RECT 394.850000 0.000000 397.550000 0.640000 ;
      RECT 391.850000 0.000000 394.550000 0.640000 ;
      RECT 388.850000 0.000000 391.550000 0.640000 ;
      RECT 385.850000 0.000000 388.550000 0.640000 ;
      RECT 382.850000 0.000000 385.550000 0.640000 ;
      RECT 379.850000 0.000000 382.550000 0.640000 ;
      RECT 376.850000 0.000000 379.550000 0.640000 ;
      RECT 373.850000 0.000000 376.550000 0.640000 ;
      RECT 370.850000 0.000000 373.550000 0.640000 ;
      RECT 367.850000 0.000000 370.550000 0.640000 ;
      RECT 364.850000 0.000000 367.550000 0.640000 ;
      RECT 361.850000 0.000000 364.550000 0.640000 ;
      RECT 358.850000 0.000000 361.550000 0.640000 ;
      RECT 355.850000 0.000000 358.550000 0.640000 ;
      RECT 352.850000 0.000000 355.550000 0.640000 ;
      RECT 349.850000 0.000000 352.550000 0.640000 ;
      RECT 346.850000 0.000000 349.550000 0.640000 ;
      RECT 343.850000 0.000000 346.550000 0.640000 ;
      RECT 340.850000 0.000000 343.550000 0.640000 ;
      RECT 337.850000 0.000000 340.550000 0.640000 ;
      RECT 334.850000 0.000000 337.550000 0.640000 ;
      RECT 331.850000 0.000000 334.550000 0.640000 ;
      RECT 328.850000 0.000000 331.550000 0.640000 ;
      RECT 325.850000 0.000000 328.550000 0.640000 ;
      RECT 322.850000 0.000000 325.550000 0.640000 ;
      RECT 319.850000 0.000000 322.550000 0.640000 ;
      RECT 316.850000 0.000000 319.550000 0.640000 ;
      RECT 313.850000 0.000000 316.550000 0.640000 ;
      RECT 310.850000 0.000000 313.550000 0.640000 ;
      RECT 307.850000 0.000000 310.550000 0.640000 ;
      RECT 304.850000 0.000000 307.550000 0.640000 ;
      RECT 301.850000 0.000000 304.550000 0.640000 ;
      RECT 298.850000 0.000000 301.550000 0.640000 ;
      RECT 295.850000 0.000000 298.550000 0.640000 ;
      RECT 292.850000 0.000000 295.550000 0.640000 ;
      RECT 289.850000 0.000000 292.550000 0.640000 ;
      RECT 286.850000 0.000000 289.550000 0.640000 ;
      RECT 283.850000 0.000000 286.550000 0.640000 ;
      RECT 280.850000 0.000000 283.550000 0.640000 ;
      RECT 277.850000 0.000000 280.550000 0.640000 ;
      RECT 274.850000 0.000000 277.550000 0.640000 ;
      RECT 271.850000 0.000000 274.550000 0.640000 ;
      RECT 268.850000 0.000000 271.550000 0.640000 ;
      RECT 265.850000 0.000000 268.550000 0.640000 ;
      RECT 262.850000 0.000000 265.550000 0.640000 ;
      RECT 259.850000 0.000000 262.550000 0.640000 ;
      RECT 256.850000 0.000000 259.550000 0.640000 ;
      RECT 253.850000 0.000000 256.550000 0.640000 ;
      RECT 250.850000 0.000000 253.550000 0.640000 ;
      RECT 247.850000 0.000000 250.550000 0.640000 ;
      RECT 244.850000 0.000000 247.550000 0.640000 ;
      RECT 241.850000 0.000000 244.550000 0.640000 ;
      RECT 238.850000 0.000000 241.550000 0.640000 ;
      RECT 235.850000 0.000000 238.550000 0.640000 ;
      RECT 232.850000 0.000000 235.550000 0.640000 ;
      RECT 229.850000 0.000000 232.550000 0.640000 ;
      RECT 226.850000 0.000000 229.550000 0.640000 ;
      RECT 223.850000 0.000000 226.550000 0.640000 ;
      RECT 220.850000 0.000000 223.550000 0.640000 ;
      RECT 217.850000 0.000000 220.550000 0.640000 ;
      RECT 214.850000 0.000000 217.550000 0.640000 ;
      RECT 211.850000 0.000000 214.550000 0.640000 ;
      RECT 208.850000 0.000000 211.550000 0.640000 ;
      RECT 205.850000 0.000000 208.550000 0.640000 ;
      RECT 202.850000 0.000000 205.550000 0.640000 ;
      RECT 199.850000 0.000000 202.550000 0.640000 ;
      RECT 196.850000 0.000000 199.550000 0.640000 ;
      RECT 193.850000 0.000000 196.550000 0.640000 ;
      RECT 190.850000 0.000000 193.550000 0.640000 ;
      RECT 187.850000 0.000000 190.550000 0.640000 ;
      RECT 184.850000 0.000000 187.550000 0.640000 ;
      RECT 181.850000 0.000000 184.550000 0.640000 ;
      RECT 178.850000 0.000000 181.550000 0.640000 ;
      RECT 175.850000 0.000000 178.550000 0.640000 ;
      RECT 172.850000 0.000000 175.550000 0.640000 ;
      RECT 169.850000 0.000000 172.550000 0.640000 ;
      RECT 166.850000 0.000000 169.550000 0.640000 ;
      RECT 163.850000 0.000000 166.550000 0.640000 ;
      RECT 160.850000 0.000000 163.550000 0.640000 ;
      RECT 157.850000 0.000000 160.550000 0.640000 ;
      RECT 154.850000 0.000000 157.550000 0.640000 ;
      RECT 151.850000 0.000000 154.550000 0.640000 ;
      RECT 148.850000 0.000000 151.550000 0.640000 ;
      RECT 145.850000 0.000000 148.550000 0.640000 ;
      RECT 142.850000 0.000000 145.550000 0.640000 ;
      RECT 139.850000 0.000000 142.550000 0.640000 ;
      RECT 136.850000 0.000000 139.550000 0.640000 ;
      RECT 133.850000 0.000000 136.550000 0.640000 ;
      RECT 130.850000 0.000000 133.550000 0.640000 ;
      RECT 0.000000 0.000000 130.550000 0.640000 ;
    LAYER M3 ;
      RECT 0.000000 420.150000 473.800000 473.600000 ;
      RECT 0.640000 419.850000 473.800000 420.150000 ;
      RECT 0.000000 415.150000 473.800000 419.850000 ;
      RECT 0.640000 414.850000 473.800000 415.150000 ;
      RECT 0.000000 410.150000 473.800000 414.850000 ;
      RECT 0.640000 409.850000 473.800000 410.150000 ;
      RECT 0.000000 405.150000 473.800000 409.850000 ;
      RECT 0.640000 404.850000 473.800000 405.150000 ;
      RECT 0.000000 400.150000 473.800000 404.850000 ;
      RECT 0.640000 399.850000 473.800000 400.150000 ;
      RECT 0.000000 395.150000 473.800000 399.850000 ;
      RECT 0.640000 394.850000 473.800000 395.150000 ;
      RECT 0.000000 390.150000 473.800000 394.850000 ;
      RECT 0.640000 389.850000 473.800000 390.150000 ;
      RECT 0.000000 385.150000 473.800000 389.850000 ;
      RECT 0.640000 384.850000 473.800000 385.150000 ;
      RECT 0.000000 380.150000 473.800000 384.850000 ;
      RECT 0.640000 379.850000 473.800000 380.150000 ;
      RECT 0.000000 375.150000 473.800000 379.850000 ;
      RECT 0.640000 374.850000 473.800000 375.150000 ;
      RECT 0.000000 370.150000 473.800000 374.850000 ;
      RECT 0.640000 369.850000 473.800000 370.150000 ;
      RECT 0.000000 365.150000 473.800000 369.850000 ;
      RECT 0.640000 364.850000 473.800000 365.150000 ;
      RECT 0.000000 360.150000 473.800000 364.850000 ;
      RECT 0.640000 359.850000 473.800000 360.150000 ;
      RECT 0.000000 355.150000 473.800000 359.850000 ;
      RECT 0.640000 354.850000 473.800000 355.150000 ;
      RECT 0.000000 350.150000 473.800000 354.850000 ;
      RECT 0.640000 349.850000 473.800000 350.150000 ;
      RECT 0.000000 345.150000 473.800000 349.850000 ;
      RECT 0.640000 344.850000 473.800000 345.150000 ;
      RECT 0.000000 340.150000 473.800000 344.850000 ;
      RECT 0.640000 339.850000 473.800000 340.150000 ;
      RECT 0.000000 335.150000 473.800000 339.850000 ;
      RECT 0.640000 334.850000 473.800000 335.150000 ;
      RECT 0.000000 330.150000 473.800000 334.850000 ;
      RECT 0.640000 329.850000 473.800000 330.150000 ;
      RECT 0.000000 325.150000 473.800000 329.850000 ;
      RECT 0.640000 324.850000 473.800000 325.150000 ;
      RECT 0.000000 320.150000 473.800000 324.850000 ;
      RECT 0.640000 319.850000 473.800000 320.150000 ;
      RECT 0.000000 315.150000 473.800000 319.850000 ;
      RECT 0.640000 314.850000 473.800000 315.150000 ;
      RECT 0.000000 310.150000 473.800000 314.850000 ;
      RECT 0.640000 309.850000 473.800000 310.150000 ;
      RECT 0.000000 305.150000 473.800000 309.850000 ;
      RECT 0.640000 304.850000 473.800000 305.150000 ;
      RECT 0.000000 300.150000 473.800000 304.850000 ;
      RECT 0.640000 299.850000 473.800000 300.150000 ;
      RECT 0.000000 295.150000 473.800000 299.850000 ;
      RECT 0.640000 294.850000 473.800000 295.150000 ;
      RECT 0.000000 290.150000 473.800000 294.850000 ;
      RECT 0.640000 289.850000 473.800000 290.150000 ;
      RECT 0.000000 285.150000 473.800000 289.850000 ;
      RECT 0.640000 284.850000 473.800000 285.150000 ;
      RECT 0.000000 280.150000 473.800000 284.850000 ;
      RECT 0.640000 279.850000 473.800000 280.150000 ;
      RECT 0.000000 275.150000 473.800000 279.850000 ;
      RECT 0.640000 274.850000 473.800000 275.150000 ;
      RECT 0.000000 270.150000 473.800000 274.850000 ;
      RECT 0.640000 269.850000 473.800000 270.150000 ;
      RECT 0.000000 265.150000 473.800000 269.850000 ;
      RECT 0.640000 264.850000 473.800000 265.150000 ;
      RECT 0.000000 260.150000 473.800000 264.850000 ;
      RECT 0.640000 259.850000 473.800000 260.150000 ;
      RECT 0.000000 255.150000 473.800000 259.850000 ;
      RECT 0.640000 254.850000 473.800000 255.150000 ;
      RECT 0.000000 250.150000 473.800000 254.850000 ;
      RECT 0.640000 249.850000 473.800000 250.150000 ;
      RECT 0.000000 245.150000 473.800000 249.850000 ;
      RECT 0.640000 244.850000 473.800000 245.150000 ;
      RECT 0.000000 240.150000 473.800000 244.850000 ;
      RECT 0.640000 239.850000 473.800000 240.150000 ;
      RECT 0.000000 235.150000 473.800000 239.850000 ;
      RECT 0.640000 234.850000 473.800000 235.150000 ;
      RECT 0.000000 230.150000 473.800000 234.850000 ;
      RECT 0.640000 229.850000 473.800000 230.150000 ;
      RECT 0.000000 225.150000 473.800000 229.850000 ;
      RECT 0.640000 224.850000 473.800000 225.150000 ;
      RECT 0.000000 220.150000 473.800000 224.850000 ;
      RECT 0.640000 219.850000 473.800000 220.150000 ;
      RECT 0.000000 215.150000 473.800000 219.850000 ;
      RECT 0.640000 214.850000 473.800000 215.150000 ;
      RECT 0.000000 210.150000 473.800000 214.850000 ;
      RECT 0.640000 209.850000 473.800000 210.150000 ;
      RECT 0.000000 205.150000 473.800000 209.850000 ;
      RECT 0.640000 204.850000 473.800000 205.150000 ;
      RECT 0.000000 200.150000 473.800000 204.850000 ;
      RECT 0.640000 199.850000 473.800000 200.150000 ;
      RECT 0.000000 195.150000 473.800000 199.850000 ;
      RECT 0.640000 194.850000 473.800000 195.150000 ;
      RECT 0.000000 190.150000 473.800000 194.850000 ;
      RECT 0.640000 189.850000 473.800000 190.150000 ;
      RECT 0.000000 185.150000 473.800000 189.850000 ;
      RECT 0.640000 184.850000 473.800000 185.150000 ;
      RECT 0.000000 180.150000 473.800000 184.850000 ;
      RECT 0.640000 179.850000 473.800000 180.150000 ;
      RECT 0.000000 175.150000 473.800000 179.850000 ;
      RECT 0.640000 174.850000 473.800000 175.150000 ;
      RECT 0.000000 170.150000 473.800000 174.850000 ;
      RECT 0.640000 169.850000 473.800000 170.150000 ;
      RECT 0.000000 165.150000 473.800000 169.850000 ;
      RECT 0.640000 164.850000 473.800000 165.150000 ;
      RECT 0.000000 160.150000 473.800000 164.850000 ;
      RECT 0.640000 159.850000 473.800000 160.150000 ;
      RECT 0.000000 155.150000 473.800000 159.850000 ;
      RECT 0.640000 154.850000 473.800000 155.150000 ;
      RECT 0.000000 150.150000 473.800000 154.850000 ;
      RECT 0.640000 149.850000 473.800000 150.150000 ;
      RECT 0.000000 145.150000 473.800000 149.850000 ;
      RECT 0.640000 144.850000 473.800000 145.150000 ;
      RECT 0.000000 140.150000 473.800000 144.850000 ;
      RECT 0.640000 139.850000 473.800000 140.150000 ;
      RECT 0.000000 135.150000 473.800000 139.850000 ;
      RECT 0.640000 134.850000 473.800000 135.150000 ;
      RECT 0.000000 130.150000 473.800000 134.850000 ;
      RECT 0.640000 129.850000 473.800000 130.150000 ;
      RECT 0.000000 125.150000 473.800000 129.850000 ;
      RECT 0.640000 124.850000 473.800000 125.150000 ;
      RECT 0.000000 120.150000 473.800000 124.850000 ;
      RECT 0.640000 119.850000 473.800000 120.150000 ;
      RECT 0.000000 115.150000 473.800000 119.850000 ;
      RECT 0.640000 114.850000 473.800000 115.150000 ;
      RECT 0.000000 110.150000 473.800000 114.850000 ;
      RECT 0.640000 109.850000 473.800000 110.150000 ;
      RECT 0.000000 105.150000 473.800000 109.850000 ;
      RECT 0.640000 104.850000 473.800000 105.150000 ;
      RECT 0.000000 100.150000 473.800000 104.850000 ;
      RECT 0.640000 99.850000 473.800000 100.150000 ;
      RECT 0.000000 95.150000 473.800000 99.850000 ;
      RECT 0.640000 94.850000 473.800000 95.150000 ;
      RECT 0.000000 90.150000 473.800000 94.850000 ;
      RECT 0.640000 89.850000 473.800000 90.150000 ;
      RECT 0.000000 85.150000 473.800000 89.850000 ;
      RECT 0.640000 84.850000 473.800000 85.150000 ;
      RECT 0.000000 80.150000 473.800000 84.850000 ;
      RECT 0.640000 79.850000 473.800000 80.150000 ;
      RECT 0.000000 75.150000 473.800000 79.850000 ;
      RECT 0.640000 74.850000 473.800000 75.150000 ;
      RECT 0.000000 70.150000 473.800000 74.850000 ;
      RECT 0.640000 69.850000 473.800000 70.150000 ;
      RECT 0.000000 65.150000 473.800000 69.850000 ;
      RECT 0.640000 64.850000 473.800000 65.150000 ;
      RECT 0.000000 60.150000 473.800000 64.850000 ;
      RECT 0.640000 59.850000 473.800000 60.150000 ;
      RECT 0.000000 55.150000 473.800000 59.850000 ;
      RECT 0.640000 54.850000 473.800000 55.150000 ;
      RECT 0.000000 50.150000 473.800000 54.850000 ;
      RECT 0.640000 49.850000 473.800000 50.150000 ;
      RECT 0.000000 45.150000 473.800000 49.850000 ;
      RECT 0.640000 44.850000 473.800000 45.150000 ;
      RECT 0.000000 40.150000 473.800000 44.850000 ;
      RECT 0.640000 39.850000 473.800000 40.150000 ;
      RECT 0.000000 35.150000 473.800000 39.850000 ;
      RECT 0.640000 34.850000 473.800000 35.150000 ;
      RECT 0.000000 30.150000 473.800000 34.850000 ;
      RECT 0.640000 29.850000 473.800000 30.150000 ;
      RECT 0.000000 25.150000 473.800000 29.850000 ;
      RECT 0.640000 24.850000 473.800000 25.150000 ;
      RECT 0.000000 20.150000 473.800000 24.850000 ;
      RECT 0.640000 19.850000 473.800000 20.150000 ;
      RECT 0.000000 15.150000 473.800000 19.850000 ;
      RECT 0.640000 14.850000 473.800000 15.150000 ;
      RECT 0.000000 10.150000 473.800000 14.850000 ;
      RECT 0.640000 9.850000 473.800000 10.150000 ;
      RECT 0.000000 0.000000 473.800000 9.850000 ;
    LAYER M4 ;
      RECT 0.000000 0.000000 473.800000 473.600000 ;
    LAYER M5 ;
      RECT 0.000000 0.000000 473.800000 473.600000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 473.800000 473.600000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 473.800000 473.600000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 473.800000 473.600000 ;
  END
END fullchip

END LIBRARY
